-- TestBench Template 

  LIBRARY ieee;
  USE ieee.std_logic_1164.ALL;
  USE ieee.numeric_std.ALL;
  use Work.My_Package.all;

  ENTITY testbench IS
  END testbench;

  ARCHITECTURE behavior OF testbench IS 

  -- Component Declaration
          COMPONENT main
			port (picture_in : in pic_type ;
					pic_out : out result_type);
          END COMPONENT;

          SIGNAL picture_in :  pic_type;
          SIGNAL pic_out :  result_type;
          
  BEGIN

  -- Component Instantiation
          uut: main PORT MAP(
                 picture_in => picture_in,
                  pic_out => pic_out
          );


  --  Test Bench Statements
     tb : PROCESS
     BEGIN
		picture_in<=((1.780000000000000000e+02,1.730000000000000000e+02,1.560000000000000000e+02,1.330000000000000000e+02,9.100000000000000000e+01,6.500000000000000000e+01,8.200000000000000000e+01,1.200000000000000000e+02,1.610000000000000000e+02,1.560000000000000000e+02,1.460000000000000000e+02,1.200000000000000000e+02,6.900000000000000000e+01,3.100000000000000000e+01,1.100000000000000000e+01,1.600000000000000000e+01,2.200000000000000000e+01,2.300000000000000000e+01,2.800000000000000000e+01,3.500000000000000000e+01,3.500000000000000000e+01,4.300000000000000000e+01,4.200000000000000000e+01,4.300000000000000000e+01,3.200000000000000000e+01,3.500000000000000000e+01,3.000000000000000000e+01,2.200000000000000000e+01,5.700000000000000000e+01,1.120000000000000000e+02,5.200000000000000000e+01,7.700000000000000000e+01,6.000000000000000000e+01,7.000000000000000000e+01,5.700000000000000000e+01,5.700000000000000000e+01,4.200000000000000000e+01,2.800000000000000000e+01,2.600000000000000000e+01,4.200000000000000000e+01,5.300000000000000000e+01,5.600000000000000000e+01,5.700000000000000000e+01,5.300000000000000000e+01,5.900000000000000000e+01,4.300000000000000000e+01,4.700000000000000000e+01,5.200000000000000000e+01,5.400000000000000000e+01,7.000000000000000000e+01,8.300000000000000000e+01,7.700000000000000000e+01,6.900000000000000000e+01,6.900000000000000000e+01,6.400000000000000000e+01,5.700000000000000000e+01,4.700000000000000000e+01,4.300000000000000000e+01,4.400000000000000000e+01,4.400000000000000000e+01,5.400000000000000000e+01,6.600000000000000000e+01,7.300000000000000000e+01,7.300000000000000000e+01,6.700000000000000000e+01,7.000000000000000000e+01,6.300000000000000000e+01,6.600000000000000000e+01,6.100000000000000000e+01,6.500000000000000000e+01,7.500000000000000000e+01,8.000000000000000000e+01,8.700000000000000000e+01,8.800000000000000000e+01,8.400000000000000000e+01,7.600000000000000000e+01,6.500000000000000000e+01,5.200000000000000000e+01,5.400000000000000000e+01,4.900000000000000000e+01,5.800000000000000000e+01,7.200000000000000000e+01,7.600000000000000000e+01,8.100000000000000000e+01,8.700000000000000000e+01,8.800000000000000000e+01,8.000000000000000000e+01,7.700000000000000000e+01,6.900000000000000000e+01,7.800000000000000000e+01,6.900000000000000000e+01,7.300000000000000000e+01,8.600000000000000000e+01,9.200000000000000000e+01,8.300000000000000000e+01,7.200000000000000000e+01,7.500000000000000000e+01,6.900000000000000000e+01,6.000000000000000000e+01,5.300000000000000000e+01,4.600000000000000000e+01,4.300000000000000000e+01,4.700000000000000000e+01,4.200000000000000000e+01,8.600000000000000000e+01,1.340000000000000000e+02,1.690000000000000000e+02,1.910000000000000000e+02,2.030000000000000000e+02,2.050000000000000000e+02,2.020000000000000000e+02,1.970000000000000000e+02,1.940000000000000000e+02,1.960000000000000000e+02,1.980000000000000000e+02,2.030000000000000000e+02,2.060000000000000000e+02,2.030000000000000000e+02,2.110000000000000000e+02,2.130000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.070000000000000000e+02,1.350000000000000000e+02,1.320000000000000000e+02,1.260000000000000000e+02),
(1.760000000000000000e+02,1.810000000000000000e+02,1.580000000000000000e+02,1.250000000000000000e+02,9.300000000000000000e+01,6.100000000000000000e+01,8.000000000000000000e+01,1.100000000000000000e+02,1.570000000000000000e+02,1.600000000000000000e+02,1.460000000000000000e+02,1.120000000000000000e+02,7.100000000000000000e+01,3.400000000000000000e+01,1.600000000000000000e+01,2.100000000000000000e+01,2.600000000000000000e+01,3.000000000000000000e+01,3.700000000000000000e+01,3.200000000000000000e+01,3.400000000000000000e+01,3.200000000000000000e+01,3.800000000000000000e+01,3.800000000000000000e+01,3.700000000000000000e+01,3.900000000000000000e+01,2.600000000000000000e+01,6.700000000000000000e+01,8.400000000000000000e+01,6.300000000000000000e+01,6.200000000000000000e+01,6.700000000000000000e+01,6.600000000000000000e+01,7.600000000000000000e+01,7.300000000000000000e+01,7.800000000000000000e+01,6.400000000000000000e+01,7.700000000000000000e+01,2.000000000000000000e+01,4.200000000000000000e+01,4.900000000000000000e+01,5.100000000000000000e+01,4.200000000000000000e+01,4.200000000000000000e+01,4.800000000000000000e+01,5.200000000000000000e+01,6.000000000000000000e+01,6.300000000000000000e+01,6.900000000000000000e+01,7.300000000000000000e+01,7.000000000000000000e+01,6.700000000000000000e+01,5.800000000000000000e+01,4.400000000000000000e+01,4.500000000000000000e+01,5.300000000000000000e+01,5.200000000000000000e+01,5.600000000000000000e+01,6.400000000000000000e+01,6.200000000000000000e+01,6.700000000000000000e+01,5.800000000000000000e+01,5.100000000000000000e+01,5.200000000000000000e+01,5.100000000000000000e+01,6.500000000000000000e+01,6.500000000000000000e+01,7.300000000000000000e+01,8.200000000000000000e+01,8.200000000000000000e+01,9.400000000000000000e+01,9.500000000000000000e+01,8.900000000000000000e+01,7.400000000000000000e+01,6.700000000000000000e+01,6.100000000000000000e+01,5.900000000000000000e+01,6.400000000000000000e+01,6.900000000000000000e+01,7.000000000000000000e+01,7.500000000000000000e+01,7.800000000000000000e+01,7.600000000000000000e+01,7.500000000000000000e+01,6.500000000000000000e+01,5.700000000000000000e+01,6.400000000000000000e+01,6.700000000000000000e+01,6.700000000000000000e+01,8.000000000000000000e+01,7.700000000000000000e+01,8.200000000000000000e+01,8.200000000000000000e+01,7.900000000000000000e+01,6.800000000000000000e+01,5.500000000000000000e+01,4.700000000000000000e+01,5.600000000000000000e+01,5.500000000000000000e+01,5.500000000000000000e+01,5.300000000000000000e+01,6.300000000000000000e+01,5.800000000000000000e+01,5.100000000000000000e+01,7.900000000000000000e+01,1.250000000000000000e+02,1.660000000000000000e+02,1.910000000000000000e+02,2.030000000000000000e+02,2.050000000000000000e+02,2.000000000000000000e+02,1.980000000000000000e+02,1.930000000000000000e+02,1.930000000000000000e+02,1.950000000000000000e+02,2.000000000000000000e+02,2.050000000000000000e+02,2.020000000000000000e+02,2.110000000000000000e+02,2.130000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.080000000000000000e+02,1.310000000000000000e+02,1.280000000000000000e+02,1.260000000000000000e+02),
(1.790000000000000000e+02,1.740000000000000000e+02,1.590000000000000000e+02,1.240000000000000000e+02,8.900000000000000000e+01,6.000000000000000000e+01,7.900000000000000000e+01,1.100000000000000000e+02,1.500000000000000000e+02,1.580000000000000000e+02,1.460000000000000000e+02,1.100000000000000000e+02,7.500000000000000000e+01,4.000000000000000000e+01,2.400000000000000000e+01,2.700000000000000000e+01,3.300000000000000000e+01,3.700000000000000000e+01,4.100000000000000000e+01,3.600000000000000000e+01,3.200000000000000000e+01,3.100000000000000000e+01,3.100000000000000000e+01,3.600000000000000000e+01,3.900000000000000000e+01,4.200000000000000000e+01,2.900000000000000000e+01,6.900000000000000000e+01,6.700000000000000000e+01,6.800000000000000000e+01,6.300000000000000000e+01,7.800000000000000000e+01,9.100000000000000000e+01,7.700000000000000000e+01,7.400000000000000000e+01,7.900000000000000000e+01,6.600000000000000000e+01,6.100000000000000000e+01,6.400000000000000000e+01,3.400000000000000000e+01,4.100000000000000000e+01,4.200000000000000000e+01,4.000000000000000000e+01,3.600000000000000000e+01,3.800000000000000000e+01,4.600000000000000000e+01,6.000000000000000000e+01,7.000000000000000000e+01,8.300000000000000000e+01,6.900000000000000000e+01,6.700000000000000000e+01,5.800000000000000000e+01,4.900000000000000000e+01,3.900000000000000000e+01,4.700000000000000000e+01,4.600000000000000000e+01,5.800000000000000000e+01,7.300000000000000000e+01,8.100000000000000000e+01,7.100000000000000000e+01,7.300000000000000000e+01,6.800000000000000000e+01,5.400000000000000000e+01,4.600000000000000000e+01,4.100000000000000000e+01,4.900000000000000000e+01,6.700000000000000000e+01,7.800000000000000000e+01,8.800000000000000000e+01,1.000000000000000000e+02,9.400000000000000000e+01,9.100000000000000000e+01,8.300000000000000000e+01,7.200000000000000000e+01,6.600000000000000000e+01,5.300000000000000000e+01,5.400000000000000000e+01,6.500000000000000000e+01,6.900000000000000000e+01,8.100000000000000000e+01,8.300000000000000000e+01,8.500000000000000000e+01,7.400000000000000000e+01,6.700000000000000000e+01,5.700000000000000000e+01,5.200000000000000000e+01,5.200000000000000000e+01,6.700000000000000000e+01,6.900000000000000000e+01,7.700000000000000000e+01,8.600000000000000000e+01,8.600000000000000000e+01,7.900000000000000000e+01,7.000000000000000000e+01,6.300000000000000000e+01,5.200000000000000000e+01,4.300000000000000000e+01,3.900000000000000000e+01,4.200000000000000000e+01,5.500000000000000000e+01,5.700000000000000000e+01,6.600000000000000000e+01,1.070000000000000000e+02,5.300000000000000000e+01,8.600000000000000000e+01,1.280000000000000000e+02,1.650000000000000000e+02,1.910000000000000000e+02,2.030000000000000000e+02,2.040000000000000000e+02,1.990000000000000000e+02,1.990000000000000000e+02,1.940000000000000000e+02,1.930000000000000000e+02,1.950000000000000000e+02,1.990000000000000000e+02,2.040000000000000000e+02,2.020000000000000000e+02,2.120000000000000000e+02,2.160000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.080000000000000000e+02,1.350000000000000000e+02,1.340000000000000000e+02,1.290000000000000000e+02),
(1.810000000000000000e+02,1.760000000000000000e+02,1.580000000000000000e+02,1.200000000000000000e+02,9.300000000000000000e+01,6.100000000000000000e+01,8.400000000000000000e+01,1.110000000000000000e+02,1.570000000000000000e+02,1.610000000000000000e+02,1.480000000000000000e+02,1.170000000000000000e+02,7.900000000000000000e+01,4.400000000000000000e+01,2.400000000000000000e+01,3.300000000000000000e+01,4.000000000000000000e+01,4.200000000000000000e+01,4.100000000000000000e+01,3.300000000000000000e+01,3.700000000000000000e+01,3.300000000000000000e+01,3.000000000000000000e+01,3.500000000000000000e+01,3.900000000000000000e+01,2.400000000000000000e+01,4.900000000000000000e+01,5.500000000000000000e+01,6.700000000000000000e+01,7.000000000000000000e+01,8.900000000000000000e+01,8.900000000000000000e+01,9.200000000000000000e+01,1.060000000000000000e+02,9.700000000000000000e+01,1.040000000000000000e+02,8.200000000000000000e+01,6.900000000000000000e+01,8.100000000000000000e+01,7.400000000000000000e+01,4.300000000000000000e+01,2.900000000000000000e+01,3.900000000000000000e+01,2.600000000000000000e+01,3.200000000000000000e+01,4.300000000000000000e+01,6.500000000000000000e+01,7.200000000000000000e+01,7.100000000000000000e+01,7.000000000000000000e+01,5.500000000000000000e+01,5.000000000000000000e+01,4.200000000000000000e+01,3.700000000000000000e+01,4.300000000000000000e+01,4.800000000000000000e+01,6.000000000000000000e+01,7.600000000000000000e+01,9.200000000000000000e+01,8.800000000000000000e+01,7.700000000000000000e+01,7.500000000000000000e+01,6.300000000000000000e+01,5.200000000000000000e+01,4.400000000000000000e+01,4.700000000000000000e+01,5.900000000000000000e+01,8.000000000000000000e+01,8.900000000000000000e+01,1.020000000000000000e+02,9.300000000000000000e+01,8.200000000000000000e+01,7.700000000000000000e+01,6.400000000000000000e+01,6.300000000000000000e+01,5.600000000000000000e+01,5.300000000000000000e+01,5.400000000000000000e+01,6.800000000000000000e+01,8.700000000000000000e+01,8.600000000000000000e+01,8.400000000000000000e+01,7.300000000000000000e+01,6.800000000000000000e+01,5.300000000000000000e+01,4.900000000000000000e+01,4.700000000000000000e+01,5.200000000000000000e+01,6.100000000000000000e+01,7.900000000000000000e+01,8.600000000000000000e+01,8.700000000000000000e+01,7.300000000000000000e+01,6.100000000000000000e+01,5.200000000000000000e+01,4.900000000000000000e+01,4.300000000000000000e+01,3.900000000000000000e+01,4.300000000000000000e+01,5.500000000000000000e+01,6.700000000000000000e+01,7.300000000000000000e+01,6.700000000000000000e+01,6.100000000000000000e+01,8.900000000000000000e+01,1.290000000000000000e+02,1.660000000000000000e+02,1.930000000000000000e+02,2.020000000000000000e+02,2.030000000000000000e+02,1.990000000000000000e+02,1.960000000000000000e+02,1.930000000000000000e+02,1.880000000000000000e+02,1.950000000000000000e+02,1.990000000000000000e+02,2.020000000000000000e+02,2.010000000000000000e+02,2.120000000000000000e+02,2.160000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.100000000000000000e+02,1.360000000000000000e+02,1.310000000000000000e+02,1.270000000000000000e+02),
(1.800000000000000000e+02,1.770000000000000000e+02,1.490000000000000000e+02,1.210000000000000000e+02,8.900000000000000000e+01,5.800000000000000000e+01,8.200000000000000000e+01,1.170000000000000000e+02,1.540000000000000000e+02,1.610000000000000000e+02,1.460000000000000000e+02,1.150000000000000000e+02,7.700000000000000000e+01,4.400000000000000000e+01,2.800000000000000000e+01,3.600000000000000000e+01,4.900000000000000000e+01,4.300000000000000000e+01,3.700000000000000000e+01,3.700000000000000000e+01,4.300000000000000000e+01,3.200000000000000000e+01,2.900000000000000000e+01,3.700000000000000000e+01,3.000000000000000000e+01,7.000000000000000000e+01,7.000000000000000000e+01,4.200000000000000000e+01,6.500000000000000000e+01,9.200000000000000000e+01,9.700000000000000000e+01,1.080000000000000000e+02,1.140000000000000000e+02,1.230000000000000000e+02,1.220000000000000000e+02,1.200000000000000000e+02,1.240000000000000000e+02,1.050000000000000000e+02,8.100000000000000000e+01,8.900000000000000000e+01,9.300000000000000000e+01,5.600000000000000000e+01,2.600000000000000000e+01,2.800000000000000000e+01,3.800000000000000000e+01,4.800000000000000000e+01,5.900000000000000000e+01,6.700000000000000000e+01,7.200000000000000000e+01,6.400000000000000000e+01,5.300000000000000000e+01,4.600000000000000000e+01,4.200000000000000000e+01,3.500000000000000000e+01,4.600000000000000000e+01,5.600000000000000000e+01,6.900000000000000000e+01,8.100000000000000000e+01,9.000000000000000000e+01,9.800000000000000000e+01,9.300000000000000000e+01,7.900000000000000000e+01,7.200000000000000000e+01,6.000000000000000000e+01,4.900000000000000000e+01,5.100000000000000000e+01,6.100000000000000000e+01,7.400000000000000000e+01,8.500000000000000000e+01,8.500000000000000000e+01,8.100000000000000000e+01,7.700000000000000000e+01,6.500000000000000000e+01,6.100000000000000000e+01,6.400000000000000000e+01,6.200000000000000000e+01,6.400000000000000000e+01,6.900000000000000000e+01,7.900000000000000000e+01,9.000000000000000000e+01,8.900000000000000000e+01,9.100000000000000000e+01,8.500000000000000000e+01,7.200000000000000000e+01,5.300000000000000000e+01,4.100000000000000000e+01,4.800000000000000000e+01,4.900000000000000000e+01,5.900000000000000000e+01,6.700000000000000000e+01,7.800000000000000000e+01,7.400000000000000000e+01,6.300000000000000000e+01,5.400000000000000000e+01,4.800000000000000000e+01,4.400000000000000000e+01,4.500000000000000000e+01,5.400000000000000000e+01,5.500000000000000000e+01,6.300000000000000000e+01,6.900000000000000000e+01,7.500000000000000000e+01,6.800000000000000000e+01,5.600000000000000000e+01,9.200000000000000000e+01,1.260000000000000000e+02,1.650000000000000000e+02,1.880000000000000000e+02,2.020000000000000000e+02,2.050000000000000000e+02,2.000000000000000000e+02,1.940000000000000000e+02,1.920000000000000000e+02,1.900000000000000000e+02,1.920000000000000000e+02,1.950000000000000000e+02,2.020000000000000000e+02,1.990000000000000000e+02,2.110000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.090000000000000000e+02,1.360000000000000000e+02,1.330000000000000000e+02,1.280000000000000000e+02),
(1.790000000000000000e+02,1.750000000000000000e+02,1.550000000000000000e+02,1.180000000000000000e+02,9.000000000000000000e+01,5.900000000000000000e+01,8.400000000000000000e+01,1.150000000000000000e+02,1.570000000000000000e+02,1.610000000000000000e+02,1.440000000000000000e+02,1.230000000000000000e+02,7.900000000000000000e+01,4.400000000000000000e+01,2.800000000000000000e+01,4.000000000000000000e+01,4.900000000000000000e+01,4.600000000000000000e+01,4.300000000000000000e+01,4.000000000000000000e+01,4.200000000000000000e+01,3.500000000000000000e+01,3.200000000000000000e+01,3.900000000000000000e+01,3.300000000000000000e+01,5.800000000000000000e+01,4.500000000000000000e+01,7.000000000000000000e+01,8.400000000000000000e+01,1.040000000000000000e+02,1.040000000000000000e+02,1.070000000000000000e+02,1.230000000000000000e+02,1.290000000000000000e+02,1.290000000000000000e+02,1.370000000000000000e+02,1.390000000000000000e+02,1.340000000000000000e+02,1.090000000000000000e+02,1.090000000000000000e+02,1.070000000000000000e+02,1.000000000000000000e+02,3.900000000000000000e+01,2.700000000000000000e+01,3.700000000000000000e+01,4.800000000000000000e+01,5.800000000000000000e+01,5.700000000000000000e+01,5.700000000000000000e+01,6.600000000000000000e+01,5.000000000000000000e+01,4.600000000000000000e+01,3.800000000000000000e+01,4.200000000000000000e+01,5.400000000000000000e+01,6.100000000000000000e+01,6.600000000000000000e+01,7.800000000000000000e+01,8.600000000000000000e+01,9.400000000000000000e+01,8.900000000000000000e+01,8.400000000000000000e+01,6.400000000000000000e+01,5.300000000000000000e+01,5.100000000000000000e+01,5.500000000000000000e+01,6.300000000000000000e+01,7.100000000000000000e+01,7.700000000000000000e+01,8.400000000000000000e+01,7.500000000000000000e+01,7.600000000000000000e+01,6.700000000000000000e+01,6.300000000000000000e+01,6.400000000000000000e+01,6.500000000000000000e+01,7.200000000000000000e+01,7.300000000000000000e+01,8.300000000000000000e+01,8.600000000000000000e+01,8.700000000000000000e+01,9.300000000000000000e+01,8.600000000000000000e+01,6.700000000000000000e+01,5.500000000000000000e+01,4.900000000000000000e+01,5.600000000000000000e+01,5.700000000000000000e+01,6.000000000000000000e+01,6.700000000000000000e+01,6.700000000000000000e+01,6.700000000000000000e+01,6.200000000000000000e+01,5.400000000000000000e+01,5.500000000000000000e+01,5.800000000000000000e+01,5.400000000000000000e+01,6.500000000000000000e+01,6.000000000000000000e+01,6.000000000000000000e+01,6.700000000000000000e+01,7.000000000000000000e+01,6.800000000000000000e+01,5.600000000000000000e+01,8.200000000000000000e+01,1.240000000000000000e+02,1.590000000000000000e+02,1.880000000000000000e+02,2.010000000000000000e+02,2.040000000000000000e+02,2.000000000000000000e+02,1.940000000000000000e+02,1.900000000000000000e+02,1.890000000000000000e+02,1.920000000000000000e+02,1.950000000000000000e+02,1.990000000000000000e+02,2.000000000000000000e+02,2.100000000000000000e+02,2.150000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.110000000000000000e+02,1.370000000000000000e+02,1.340000000000000000e+02,1.300000000000000000e+02),
(1.820000000000000000e+02,1.680000000000000000e+02,1.570000000000000000e+02,1.190000000000000000e+02,8.700000000000000000e+01,5.800000000000000000e+01,8.400000000000000000e+01,1.140000000000000000e+02,1.550000000000000000e+02,1.610000000000000000e+02,1.430000000000000000e+02,1.130000000000000000e+02,7.900000000000000000e+01,4.200000000000000000e+01,2.500000000000000000e+01,3.200000000000000000e+01,3.700000000000000000e+01,4.200000000000000000e+01,4.400000000000000000e+01,4.400000000000000000e+01,4.100000000000000000e+01,3.500000000000000000e+01,3.700000000000000000e+01,3.500000000000000000e+01,7.600000000000000000e+01,7.800000000000000000e+01,5.100000000000000000e+01,7.300000000000000000e+01,9.100000000000000000e+01,1.070000000000000000e+02,1.160000000000000000e+02,1.200000000000000000e+02,1.270000000000000000e+02,1.320000000000000000e+02,1.280000000000000000e+02,1.490000000000000000e+02,1.390000000000000000e+02,1.320000000000000000e+02,1.190000000000000000e+02,1.260000000000000000e+02,8.700000000000000000e+01,1.000000000000000000e+02,9.900000000000000000e+01,2.700000000000000000e+01,4.700000000000000000e+01,5.100000000000000000e+01,4.700000000000000000e+01,4.300000000000000000e+01,4.000000000000000000e+01,4.200000000000000000e+01,4.600000000000000000e+01,5.200000000000000000e+01,5.600000000000000000e+01,6.400000000000000000e+01,6.400000000000000000e+01,6.700000000000000000e+01,6.000000000000000000e+01,5.400000000000000000e+01,6.300000000000000000e+01,8.000000000000000000e+01,8.500000000000000000e+01,8.300000000000000000e+01,7.700000000000000000e+01,6.200000000000000000e+01,5.700000000000000000e+01,5.700000000000000000e+01,6.200000000000000000e+01,5.900000000000000000e+01,6.100000000000000000e+01,6.000000000000000000e+01,6.100000000000000000e+01,7.100000000000000000e+01,6.600000000000000000e+01,6.500000000000000000e+01,8.000000000000000000e+01,7.400000000000000000e+01,7.900000000000000000e+01,6.900000000000000000e+01,7.600000000000000000e+01,7.100000000000000000e+01,7.200000000000000000e+01,7.500000000000000000e+01,8.500000000000000000e+01,7.400000000000000000e+01,6.900000000000000000e+01,6.400000000000000000e+01,6.300000000000000000e+01,6.200000000000000000e+01,5.600000000000000000e+01,5.900000000000000000e+01,5.500000000000000000e+01,5.100000000000000000e+01,5.400000000000000000e+01,6.100000000000000000e+01,6.200000000000000000e+01,7.600000000000000000e+01,7.700000000000000000e+01,8.000000000000000000e+01,6.800000000000000000e+01,6.300000000000000000e+01,5.600000000000000000e+01,4.700000000000000000e+01,5.600000000000000000e+01,4.900000000000000000e+01,8.000000000000000000e+01,1.190000000000000000e+02,1.580000000000000000e+02,1.870000000000000000e+02,1.940000000000000000e+02,1.990000000000000000e+02,2.000000000000000000e+02,1.920000000000000000e+02,1.880000000000000000e+02,1.860000000000000000e+02,1.830000000000000000e+02,1.880000000000000000e+02,1.930000000000000000e+02,1.960000000000000000e+02,2.080000000000000000e+02,2.150000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.100000000000000000e+02,1.390000000000000000e+02,1.370000000000000000e+02,1.300000000000000000e+02),
(1.770000000000000000e+02,1.700000000000000000e+02,1.540000000000000000e+02,1.190000000000000000e+02,8.900000000000000000e+01,5.600000000000000000e+01,8.300000000000000000e+01,1.140000000000000000e+02,1.570000000000000000e+02,1.590000000000000000e+02,1.510000000000000000e+02,1.110000000000000000e+02,7.300000000000000000e+01,3.900000000000000000e+01,2.000000000000000000e+01,2.200000000000000000e+01,3.200000000000000000e+01,3.600000000000000000e+01,3.800000000000000000e+01,4.100000000000000000e+01,4.400000000000000000e+01,4.400000000000000000e+01,4.200000000000000000e+01,3.200000000000000000e+01,1.060000000000000000e+02,6.300000000000000000e+01,7.900000000000000000e+01,9.000000000000000000e+01,9.800000000000000000e+01,1.030000000000000000e+02,1.200000000000000000e+02,1.340000000000000000e+02,1.320000000000000000e+02,1.320000000000000000e+02,1.410000000000000000e+02,1.410000000000000000e+02,1.320000000000000000e+02,1.310000000000000000e+02,1.250000000000000000e+02,1.340000000000000000e+02,1.040000000000000000e+02,1.130000000000000000e+02,1.160000000000000000e+02,7.500000000000000000e+01,3.800000000000000000e+01,4.500000000000000000e+01,4.600000000000000000e+01,4.100000000000000000e+01,3.300000000000000000e+01,3.700000000000000000e+01,4.300000000000000000e+01,6.200000000000000000e+01,6.400000000000000000e+01,7.300000000000000000e+01,6.800000000000000000e+01,5.900000000000000000e+01,5.600000000000000000e+01,4.100000000000000000e+01,4.600000000000000000e+01,6.700000000000000000e+01,6.300000000000000000e+01,7.700000000000000000e+01,8.300000000000000000e+01,7.700000000000000000e+01,7.100000000000000000e+01,5.600000000000000000e+01,5.800000000000000000e+01,6.000000000000000000e+01,4.500000000000000000e+01,4.700000000000000000e+01,5.300000000000000000e+01,6.100000000000000000e+01,7.400000000000000000e+01,8.800000000000000000e+01,9.900000000000000000e+01,9.700000000000000000e+01,8.600000000000000000e+01,6.800000000000000000e+01,5.900000000000000000e+01,5.800000000000000000e+01,5.500000000000000000e+01,6.300000000000000000e+01,7.600000000000000000e+01,7.700000000000000000e+01,7.700000000000000000e+01,7.900000000000000000e+01,6.700000000000000000e+01,5.700000000000000000e+01,5.400000000000000000e+01,4.600000000000000000e+01,4.200000000000000000e+01,4.400000000000000000e+01,5.200000000000000000e+01,6.000000000000000000e+01,7.800000000000000000e+01,9.000000000000000000e+01,8.900000000000000000e+01,7.700000000000000000e+01,7.500000000000000000e+01,6.200000000000000000e+01,4.900000000000000000e+01,3.400000000000000000e+01,4.300000000000000000e+01,3.900000000000000000e+01,6.800000000000000000e+01,1.080000000000000000e+02,1.350000000000000000e+02,1.410000000000000000e+02,1.590000000000000000e+02,1.760000000000000000e+02,1.750000000000000000e+02,1.660000000000000000e+02,1.540000000000000000e+02,1.490000000000000000e+02,1.590000000000000000e+02,1.780000000000000000e+02,1.880000000000000000e+02,1.900000000000000000e+02,2.050000000000000000e+02,2.150000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.120000000000000000e+02,1.440000000000000000e+02,1.320000000000000000e+02,1.290000000000000000e+02),
(1.760000000000000000e+02,1.700000000000000000e+02,1.470000000000000000e+02,1.110000000000000000e+02,8.500000000000000000e+01,5.700000000000000000e+01,7.800000000000000000e+01,1.130000000000000000e+02,1.520000000000000000e+02,1.600000000000000000e+02,1.450000000000000000e+02,1.110000000000000000e+02,6.600000000000000000e+01,3.100000000000000000e+01,1.400000000000000000e+01,2.000000000000000000e+01,2.300000000000000000e+01,2.600000000000000000e+01,3.400000000000000000e+01,4.000000000000000000e+01,4.300000000000000000e+01,5.300000000000000000e+01,5.100000000000000000e+01,5.000000000000000000e+01,9.200000000000000000e+01,4.600000000000000000e+01,8.800000000000000000e+01,8.900000000000000000e+01,1.000000000000000000e+02,1.150000000000000000e+02,1.230000000000000000e+02,1.390000000000000000e+02,1.420000000000000000e+02,1.530000000000000000e+02,1.500000000000000000e+02,1.570000000000000000e+02,1.560000000000000000e+02,1.320000000000000000e+02,1.440000000000000000e+02,1.380000000000000000e+02,1.030000000000000000e+02,1.160000000000000000e+02,1.010000000000000000e+02,1.230000000000000000e+02,6.400000000000000000e+01,3.900000000000000000e+01,4.400000000000000000e+01,4.500000000000000000e+01,3.100000000000000000e+01,3.600000000000000000e+01,3.800000000000000000e+01,5.800000000000000000e+01,7.000000000000000000e+01,7.000000000000000000e+01,6.400000000000000000e+01,5.500000000000000000e+01,4.500000000000000000e+01,4.300000000000000000e+01,4.400000000000000000e+01,5.300000000000000000e+01,5.500000000000000000e+01,6.100000000000000000e+01,7.800000000000000000e+01,8.000000000000000000e+01,7.400000000000000000e+01,5.200000000000000000e+01,4.800000000000000000e+01,4.700000000000000000e+01,4.300000000000000000e+01,4.000000000000000000e+01,4.300000000000000000e+01,5.300000000000000000e+01,5.700000000000000000e+01,8.200000000000000000e+01,1.020000000000000000e+02,9.300000000000000000e+01,7.500000000000000000e+01,6.000000000000000000e+01,4.700000000000000000e+01,5.000000000000000000e+01,4.400000000000000000e+01,5.500000000000000000e+01,6.800000000000000000e+01,8.000000000000000000e+01,8.300000000000000000e+01,7.900000000000000000e+01,6.700000000000000000e+01,5.500000000000000000e+01,4.700000000000000000e+01,4.000000000000000000e+01,3.600000000000000000e+01,4.300000000000000000e+01,4.600000000000000000e+01,6.500000000000000000e+01,7.500000000000000000e+01,9.300000000000000000e+01,8.800000000000000000e+01,7.300000000000000000e+01,6.500000000000000000e+01,5.200000000000000000e+01,3.900000000000000000e+01,3.400000000000000000e+01,3.200000000000000000e+01,3.200000000000000000e+01,5.300000000000000000e+01,9.200000000000000000e+01,9.300000000000000000e+01,1.030000000000000000e+02,1.160000000000000000e+02,1.220000000000000000e+02,1.110000000000000000e+02,9.100000000000000000e+01,9.400000000000000000e+01,1.230000000000000000e+02,1.550000000000000000e+02,1.770000000000000000e+02,1.920000000000000000e+02,1.920000000000000000e+02,2.050000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.150000000000000000e+02,2.130000000000000000e+02,2.120000000000000000e+02,1.350000000000000000e+02,1.330000000000000000e+02,1.350000000000000000e+02),
(1.780000000000000000e+02,1.690000000000000000e+02,1.490000000000000000e+02,1.090000000000000000e+02,8.100000000000000000e+01,5.500000000000000000e+01,8.500000000000000000e+01,1.080000000000000000e+02,1.510000000000000000e+02,1.550000000000000000e+02,1.450000000000000000e+02,1.120000000000000000e+02,6.500000000000000000e+01,3.000000000000000000e+01,1.800000000000000000e+01,1.700000000000000000e+01,2.100000000000000000e+01,2.400000000000000000e+01,2.600000000000000000e+01,3.700000000000000000e+01,4.300000000000000000e+01,5.600000000000000000e+01,4.500000000000000000e+01,9.500000000000000000e+01,7.600000000000000000e+01,7.600000000000000000e+01,1.010000000000000000e+02,1.080000000000000000e+02,1.210000000000000000e+02,1.240000000000000000e+02,1.310000000000000000e+02,1.440000000000000000e+02,1.350000000000000000e+02,1.400000000000000000e+02,1.580000000000000000e+02,1.450000000000000000e+02,1.510000000000000000e+02,1.490000000000000000e+02,1.450000000000000000e+02,1.530000000000000000e+02,1.480000000000000000e+02,1.380000000000000000e+02,1.080000000000000000e+02,1.160000000000000000e+02,8.300000000000000000e+01,5.500000000000000000e+01,4.200000000000000000e+01,4.000000000000000000e+01,3.300000000000000000e+01,3.300000000000000000e+01,4.300000000000000000e+01,6.000000000000000000e+01,6.300000000000000000e+01,7.500000000000000000e+01,6.600000000000000000e+01,5.400000000000000000e+01,4.500000000000000000e+01,3.800000000000000000e+01,3.900000000000000000e+01,4.900000000000000000e+01,5.300000000000000000e+01,5.900000000000000000e+01,7.200000000000000000e+01,7.200000000000000000e+01,7.200000000000000000e+01,5.200000000000000000e+01,4.500000000000000000e+01,3.800000000000000000e+01,2.900000000000000000e+01,3.300000000000000000e+01,3.800000000000000000e+01,4.300000000000000000e+01,6.000000000000000000e+01,7.600000000000000000e+01,9.200000000000000000e+01,8.300000000000000000e+01,6.900000000000000000e+01,4.900000000000000000e+01,4.100000000000000000e+01,4.400000000000000000e+01,3.700000000000000000e+01,4.400000000000000000e+01,5.300000000000000000e+01,7.400000000000000000e+01,7.600000000000000000e+01,7.300000000000000000e+01,6.700000000000000000e+01,5.200000000000000000e+01,4.900000000000000000e+01,3.600000000000000000e+01,3.400000000000000000e+01,3.900000000000000000e+01,4.700000000000000000e+01,5.900000000000000000e+01,7.200000000000000000e+01,8.400000000000000000e+01,8.300000000000000000e+01,7.200000000000000000e+01,6.100000000000000000e+01,4.700000000000000000e+01,3.700000000000000000e+01,2.400000000000000000e+01,3.800000000000000000e+01,5.200000000000000000e+01,7.800000000000000000e+01,8.700000000000000000e+01,8.400000000000000000e+01,1.030000000000000000e+02,8.600000000000000000e+01,1.040000000000000000e+02,1.100000000000000000e+02,9.800000000000000000e+01,8.400000000000000000e+01,1.340000000000000000e+02,1.700000000000000000e+02,1.850000000000000000e+02,1.930000000000000000e+02,1.910000000000000000e+02,2.020000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.150000000000000000e+02,2.130000000000000000e+02,2.120000000000000000e+02,1.290000000000000000e+02,1.350000000000000000e+02,1.300000000000000000e+02),
(1.740000000000000000e+02,1.700000000000000000e+02,1.450000000000000000e+02,1.020000000000000000e+02,8.100000000000000000e+01,5.200000000000000000e+01,7.900000000000000000e+01,1.160000000000000000e+02,1.530000000000000000e+02,1.550000000000000000e+02,1.460000000000000000e+02,1.130000000000000000e+02,6.900000000000000000e+01,2.400000000000000000e+01,1.100000000000000000e+01,1.600000000000000000e+01,2.100000000000000000e+01,2.400000000000000000e+01,2.600000000000000000e+01,3.800000000000000000e+01,4.300000000000000000e+01,4.700000000000000000e+01,4.500000000000000000e+01,1.070000000000000000e+02,6.200000000000000000e+01,8.800000000000000000e+01,1.090000000000000000e+02,1.130000000000000000e+02,1.320000000000000000e+02,1.340000000000000000e+02,1.330000000000000000e+02,1.480000000000000000e+02,1.450000000000000000e+02,1.440000000000000000e+02,1.470000000000000000e+02,1.490000000000000000e+02,1.440000000000000000e+02,1.520000000000000000e+02,1.490000000000000000e+02,1.530000000000000000e+02,1.500000000000000000e+02,1.480000000000000000e+02,1.460000000000000000e+02,8.400000000000000000e+01,1.050000000000000000e+02,9.200000000000000000e+01,4.100000000000000000e+01,3.100000000000000000e+01,2.900000000000000000e+01,3.500000000000000000e+01,4.300000000000000000e+01,5.000000000000000000e+01,6.300000000000000000e+01,6.800000000000000000e+01,6.400000000000000000e+01,5.500000000000000000e+01,4.600000000000000000e+01,3.400000000000000000e+01,3.900000000000000000e+01,5.200000000000000000e+01,5.500000000000000000e+01,6.300000000000000000e+01,7.000000000000000000e+01,6.700000000000000000e+01,6.200000000000000000e+01,5.900000000000000000e+01,4.400000000000000000e+01,3.300000000000000000e+01,2.600000000000000000e+01,2.900000000000000000e+01,3.600000000000000000e+01,4.600000000000000000e+01,6.100000000000000000e+01,6.900000000000000000e+01,7.700000000000000000e+01,8.000000000000000000e+01,7.100000000000000000e+01,5.300000000000000000e+01,4.200000000000000000e+01,4.100000000000000000e+01,3.900000000000000000e+01,4.700000000000000000e+01,6.500000000000000000e+01,7.200000000000000000e+01,8.000000000000000000e+01,7.100000000000000000e+01,7.100000000000000000e+01,5.700000000000000000e+01,4.700000000000000000e+01,3.300000000000000000e+01,3.100000000000000000e+01,3.400000000000000000e+01,5.300000000000000000e+01,6.000000000000000000e+01,7.200000000000000000e+01,7.700000000000000000e+01,7.900000000000000000e+01,7.300000000000000000e+01,5.800000000000000000e+01,4.700000000000000000e+01,4.100000000000000000e+01,6.900000000000000000e+01,1.060000000000000000e+02,1.170000000000000000e+02,1.000000000000000000e+02,1.020000000000000000e+02,1.010000000000000000e+02,8.800000000000000000e+01,8.700000000000000000e+01,7.600000000000000000e+01,9.200000000000000000e+01,9.800000000000000000e+01,9.700000000000000000e+01,1.560000000000000000e+02,1.790000000000000000e+02,1.850000000000000000e+02,1.910000000000000000e+02,1.880000000000000000e+02,1.980000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.120000000000000000e+02,2.120000000000000000e+02,1.280000000000000000e+02,1.320000000000000000e+02,1.470000000000000000e+02),
(1.720000000000000000e+02,1.670000000000000000e+02,1.420000000000000000e+02,1.030000000000000000e+02,7.800000000000000000e+01,4.800000000000000000e+01,7.500000000000000000e+01,1.050000000000000000e+02,1.490000000000000000e+02,1.580000000000000000e+02,1.440000000000000000e+02,1.100000000000000000e+02,6.300000000000000000e+01,3.600000000000000000e+01,1.100000000000000000e+01,2.600000000000000000e+01,2.100000000000000000e+01,2.700000000000000000e+01,2.900000000000000000e+01,3.500000000000000000e+01,3.800000000000000000e+01,3.700000000000000000e+01,4.300000000000000000e+01,9.100000000000000000e+01,7.800000000000000000e+01,9.900000000000000000e+01,1.080000000000000000e+02,1.130000000000000000e+02,1.250000000000000000e+02,1.370000000000000000e+02,1.410000000000000000e+02,1.460000000000000000e+02,1.620000000000000000e+02,1.660000000000000000e+02,1.600000000000000000e+02,1.600000000000000000e+02,1.620000000000000000e+02,1.570000000000000000e+02,1.630000000000000000e+02,1.600000000000000000e+02,1.580000000000000000e+02,1.670000000000000000e+02,1.480000000000000000e+02,8.900000000000000000e+01,8.700000000000000000e+01,1.110000000000000000e+02,4.600000000000000000e+01,3.500000000000000000e+01,3.700000000000000000e+01,3.900000000000000000e+01,4.200000000000000000e+01,4.200000000000000000e+01,5.000000000000000000e+01,4.700000000000000000e+01,5.100000000000000000e+01,4.500000000000000000e+01,4.300000000000000000e+01,4.000000000000000000e+01,4.400000000000000000e+01,5.000000000000000000e+01,5.900000000000000000e+01,5.900000000000000000e+01,6.000000000000000000e+01,4.800000000000000000e+01,4.700000000000000000e+01,4.500000000000000000e+01,3.900000000000000000e+01,2.900000000000000000e+01,3.100000000000000000e+01,3.400000000000000000e+01,4.100000000000000000e+01,4.300000000000000000e+01,5.800000000000000000e+01,6.300000000000000000e+01,6.500000000000000000e+01,6.200000000000000000e+01,6.000000000000000000e+01,4.600000000000000000e+01,3.900000000000000000e+01,4.100000000000000000e+01,3.800000000000000000e+01,5.300000000000000000e+01,5.800000000000000000e+01,6.500000000000000000e+01,6.100000000000000000e+01,5.800000000000000000e+01,5.200000000000000000e+01,5.200000000000000000e+01,4.400000000000000000e+01,3.600000000000000000e+01,3.100000000000000000e+01,4.000000000000000000e+01,5.300000000000000000e+01,5.800000000000000000e+01,5.500000000000000000e+01,5.300000000000000000e+01,5.600000000000000000e+01,5.200000000000000000e+01,6.000000000000000000e+01,8.300000000000000000e+01,1.030000000000000000e+02,1.220000000000000000e+02,1.280000000000000000e+02,1.380000000000000000e+02,1.440000000000000000e+02,1.420000000000000000e+02,1.200000000000000000e+02,1.030000000000000000e+02,9.200000000000000000e+01,8.500000000000000000e+01,7.800000000000000000e+01,8.500000000000000000e+01,9.100000000000000000e+01,1.560000000000000000e+02,1.770000000000000000e+02,1.840000000000000000e+02,1.870000000000000000e+02,1.870000000000000000e+02,1.940000000000000000e+02,2.150000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.120000000000000000e+02,2.110000000000000000e+02,1.310000000000000000e+02,1.310000000000000000e+02,1.270000000000000000e+02),
(1.690000000000000000e+02,1.630000000000000000e+02,1.390000000000000000e+02,1.000000000000000000e+02,7.400000000000000000e+01,5.100000000000000000e+01,8.200000000000000000e+01,1.130000000000000000e+02,1.510000000000000000e+02,1.580000000000000000e+02,1.430000000000000000e+02,1.130000000000000000e+02,6.700000000000000000e+01,3.200000000000000000e+01,1.700000000000000000e+01,2.200000000000000000e+01,2.400000000000000000e+01,2.600000000000000000e+01,3.000000000000000000e+01,3.100000000000000000e+01,3.000000000000000000e+01,2.600000000000000000e+01,5.900000000000000000e+01,7.200000000000000000e+01,8.200000000000000000e+01,9.100000000000000000e+01,1.070000000000000000e+02,1.070000000000000000e+02,1.220000000000000000e+02,1.430000000000000000e+02,1.530000000000000000e+02,1.540000000000000000e+02,1.650000000000000000e+02,1.690000000000000000e+02,1.600000000000000000e+02,1.560000000000000000e+02,1.550000000000000000e+02,1.450000000000000000e+02,1.540000000000000000e+02,1.580000000000000000e+02,1.530000000000000000e+02,1.420000000000000000e+02,1.450000000000000000e+02,1.170000000000000000e+02,8.400000000000000000e+01,1.260000000000000000e+02,9.500000000000000000e+01,5.600000000000000000e+01,4.500000000000000000e+01,4.300000000000000000e+01,3.900000000000000000e+01,3.300000000000000000e+01,3.100000000000000000e+01,2.800000000000000000e+01,4.000000000000000000e+01,4.000000000000000000e+01,4.100000000000000000e+01,5.400000000000000000e+01,5.500000000000000000e+01,5.300000000000000000e+01,5.600000000000000000e+01,5.400000000000000000e+01,3.800000000000000000e+01,3.000000000000000000e+01,2.800000000000000000e+01,3.700000000000000000e+01,3.800000000000000000e+01,4.100000000000000000e+01,4.400000000000000000e+01,4.500000000000000000e+01,3.800000000000000000e+01,4.400000000000000000e+01,4.300000000000000000e+01,4.200000000000000000e+01,4.200000000000000000e+01,4.100000000000000000e+01,4.600000000000000000e+01,4.200000000000000000e+01,4.700000000000000000e+01,5.400000000000000000e+01,5.100000000000000000e+01,5.300000000000000000e+01,5.200000000000000000e+01,5.300000000000000000e+01,4.300000000000000000e+01,3.400000000000000000e+01,4.100000000000000000e+01,3.900000000000000000e+01,3.800000000000000000e+01,4.000000000000000000e+01,4.400000000000000000e+01,4.600000000000000000e+01,4.900000000000000000e+01,4.800000000000000000e+01,4.400000000000000000e+01,3.800000000000000000e+01,4.500000000000000000e+01,6.800000000000000000e+01,1.230000000000000000e+02,1.260000000000000000e+02,1.310000000000000000e+02,1.530000000000000000e+02,1.640000000000000000e+02,1.650000000000000000e+02,1.460000000000000000e+02,1.270000000000000000e+02,1.260000000000000000e+02,1.160000000000000000e+02,1.120000000000000000e+02,9.600000000000000000e+01,9.300000000000000000e+01,9.000000000000000000e+01,9.800000000000000000e+01,1.700000000000000000e+02,1.750000000000000000e+02,1.830000000000000000e+02,1.870000000000000000e+02,1.820000000000000000e+02,1.900000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.100000000000000000e+02,1.270000000000000000e+02,1.250000000000000000e+02,1.220000000000000000e+02),
(1.700000000000000000e+02,1.590000000000000000e+02,1.350000000000000000e+02,9.800000000000000000e+01,7.300000000000000000e+01,5.200000000000000000e+01,7.900000000000000000e+01,1.160000000000000000e+02,1.560000000000000000e+02,1.540000000000000000e+02,1.460000000000000000e+02,1.120000000000000000e+02,6.900000000000000000e+01,3.900000000000000000e+01,1.900000000000000000e+01,2.600000000000000000e+01,3.600000000000000000e+01,3.500000000000000000e+01,2.800000000000000000e+01,3.200000000000000000e+01,2.300000000000000000e+01,2.400000000000000000e+01,8.200000000000000000e+01,7.200000000000000000e+01,1.060000000000000000e+02,1.140000000000000000e+02,1.040000000000000000e+02,1.060000000000000000e+02,1.250000000000000000e+02,1.440000000000000000e+02,1.510000000000000000e+02,1.500000000000000000e+02,1.760000000000000000e+02,1.750000000000000000e+02,1.850000000000000000e+02,1.790000000000000000e+02,1.660000000000000000e+02,1.670000000000000000e+02,1.580000000000000000e+02,1.640000000000000000e+02,1.550000000000000000e+02,1.480000000000000000e+02,1.610000000000000000e+02,1.480000000000000000e+02,1.060000000000000000e+02,1.080000000000000000e+02,1.240000000000000000e+02,6.300000000000000000e+01,5.000000000000000000e+01,4.700000000000000000e+01,3.000000000000000000e+01,2.700000000000000000e+01,3.200000000000000000e+01,2.700000000000000000e+01,3.200000000000000000e+01,3.600000000000000000e+01,4.600000000000000000e+01,5.400000000000000000e+01,6.600000000000000000e+01,6.200000000000000000e+01,5.500000000000000000e+01,4.600000000000000000e+01,3.600000000000000000e+01,3.200000000000000000e+01,2.600000000000000000e+01,2.900000000000000000e+01,3.200000000000000000e+01,4.100000000000000000e+01,4.500000000000000000e+01,5.000000000000000000e+01,4.000000000000000000e+01,4.700000000000000000e+01,3.700000000000000000e+01,3.500000000000000000e+01,3.800000000000000000e+01,4.000000000000000000e+01,3.400000000000000000e+01,3.900000000000000000e+01,5.200000000000000000e+01,6.200000000000000000e+01,6.400000000000000000e+01,5.400000000000000000e+01,4.900000000000000000e+01,4.400000000000000000e+01,4.000000000000000000e+01,3.100000000000000000e+01,3.200000000000000000e+01,3.100000000000000000e+01,3.300000000000000000e+01,4.100000000000000000e+01,5.100000000000000000e+01,5.100000000000000000e+01,4.300000000000000000e+01,4.200000000000000000e+01,4.300000000000000000e+01,4.500000000000000000e+01,9.700000000000000000e+01,1.100000000000000000e+02,1.250000000000000000e+02,1.320000000000000000e+02,1.640000000000000000e+02,1.770000000000000000e+02,1.530000000000000000e+02,1.350000000000000000e+02,1.300000000000000000e+02,1.050000000000000000e+02,9.700000000000000000e+01,1.100000000000000000e+02,1.090000000000000000e+02,1.100000000000000000e+02,1.090000000000000000e+02,1.060000000000000000e+02,1.190000000000000000e+02,1.700000000000000000e+02,1.770000000000000000e+02,1.810000000000000000e+02,1.860000000000000000e+02,1.890000000000000000e+02,1.900000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.110000000000000000e+02,1.260000000000000000e+02,1.250000000000000000e+02,1.250000000000000000e+02),
(1.710000000000000000e+02,1.630000000000000000e+02,1.290000000000000000e+02,9.300000000000000000e+01,7.100000000000000000e+01,5.500000000000000000e+01,7.800000000000000000e+01,1.050000000000000000e+02,1.540000000000000000e+02,1.600000000000000000e+02,1.470000000000000000e+02,1.140000000000000000e+02,7.000000000000000000e+01,3.800000000000000000e+01,1.800000000000000000e+01,2.700000000000000000e+01,3.600000000000000000e+01,2.900000000000000000e+01,2.500000000000000000e+01,2.400000000000000000e+01,2.300000000000000000e+01,2.700000000000000000e+01,8.200000000000000000e+01,7.900000000000000000e+01,1.080000000000000000e+02,1.080000000000000000e+02,1.090000000000000000e+02,1.150000000000000000e+02,1.220000000000000000e+02,1.300000000000000000e+02,1.560000000000000000e+02,1.830000000000000000e+02,1.770000000000000000e+02,1.620000000000000000e+02,1.680000000000000000e+02,1.710000000000000000e+02,1.770000000000000000e+02,1.820000000000000000e+02,1.790000000000000000e+02,1.830000000000000000e+02,1.680000000000000000e+02,1.490000000000000000e+02,1.430000000000000000e+02,1.340000000000000000e+02,1.560000000000000000e+02,1.260000000000000000e+02,1.210000000000000000e+02,1.090000000000000000e+02,4.500000000000000000e+01,4.600000000000000000e+01,2.600000000000000000e+01,2.500000000000000000e+01,2.800000000000000000e+01,2.500000000000000000e+01,2.700000000000000000e+01,3.000000000000000000e+01,3.600000000000000000e+01,4.500000000000000000e+01,5.700000000000000000e+01,5.500000000000000000e+01,4.200000000000000000e+01,3.600000000000000000e+01,3.200000000000000000e+01,3.000000000000000000e+01,2.300000000000000000e+01,2.500000000000000000e+01,3.000000000000000000e+01,4.100000000000000000e+01,4.800000000000000000e+01,4.700000000000000000e+01,4.600000000000000000e+01,3.600000000000000000e+01,3.400000000000000000e+01,3.400000000000000000e+01,3.600000000000000000e+01,2.600000000000000000e+01,2.700000000000000000e+01,3.100000000000000000e+01,4.100000000000000000e+01,5.900000000000000000e+01,6.000000000000000000e+01,4.900000000000000000e+01,4.300000000000000000e+01,4.400000000000000000e+01,4.100000000000000000e+01,3.000000000000000000e+01,2.800000000000000000e+01,2.700000000000000000e+01,3.000000000000000000e+01,4.200000000000000000e+01,5.600000000000000000e+01,5.100000000000000000e+01,4.300000000000000000e+01,3.700000000000000000e+01,6.100000000000000000e+01,1.240000000000000000e+02,1.470000000000000000e+02,1.160000000000000000e+02,1.160000000000000000e+02,1.600000000000000000e+02,1.670000000000000000e+02,1.580000000000000000e+02,1.430000000000000000e+02,1.360000000000000000e+02,1.190000000000000000e+02,1.260000000000000000e+02,1.250000000000000000e+02,1.230000000000000000e+02,1.140000000000000000e+02,1.110000000000000000e+02,1.210000000000000000e+02,1.110000000000000000e+02,1.220000000000000000e+02,1.720000000000000000e+02,1.770000000000000000e+02,1.800000000000000000e+02,1.850000000000000000e+02,1.880000000000000000e+02,1.860000000000000000e+02,2.120000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.120000000000000000e+02,1.870000000000000000e+02,1.850000000000000000e+02,1.850000000000000000e+02),
(1.720000000000000000e+02,1.600000000000000000e+02,1.360000000000000000e+02,9.200000000000000000e+01,7.500000000000000000e+01,5.500000000000000000e+01,7.800000000000000000e+01,1.110000000000000000e+02,1.570000000000000000e+02,1.600000000000000000e+02,1.470000000000000000e+02,1.110000000000000000e+02,7.000000000000000000e+01,3.500000000000000000e+01,2.100000000000000000e+01,2.700000000000000000e+01,3.400000000000000000e+01,2.900000000000000000e+01,3.000000000000000000e+01,2.900000000000000000e+01,2.000000000000000000e+01,7.800000000000000000e+01,7.700000000000000000e+01,9.600000000000000000e+01,1.060000000000000000e+02,9.500000000000000000e+01,1.020000000000000000e+02,1.280000000000000000e+02,1.410000000000000000e+02,1.550000000000000000e+02,1.610000000000000000e+02,1.840000000000000000e+02,2.000000000000000000e+02,2.010000000000000000e+02,1.900000000000000000e+02,1.880000000000000000e+02,1.890000000000000000e+02,1.900000000000000000e+02,1.890000000000000000e+02,1.820000000000000000e+02,1.800000000000000000e+02,1.730000000000000000e+02,1.490000000000000000e+02,1.190000000000000000e+02,1.320000000000000000e+02,1.390000000000000000e+02,1.180000000000000000e+02,1.370000000000000000e+02,6.900000000000000000e+01,3.400000000000000000e+01,4.100000000000000000e+01,3.100000000000000000e+01,2.700000000000000000e+01,2.100000000000000000e+01,2.700000000000000000e+01,3.600000000000000000e+01,4.200000000000000000e+01,4.200000000000000000e+01,5.900000000000000000e+01,4.800000000000000000e+01,4.500000000000000000e+01,3.600000000000000000e+01,2.900000000000000000e+01,2.400000000000000000e+01,2.000000000000000000e+01,2.500000000000000000e+01,3.200000000000000000e+01,4.200000000000000000e+01,4.500000000000000000e+01,5.200000000000000000e+01,4.100000000000000000e+01,3.900000000000000000e+01,3.800000000000000000e+01,2.900000000000000000e+01,2.800000000000000000e+01,2.600000000000000000e+01,3.300000000000000000e+01,3.400000000000000000e+01,4.000000000000000000e+01,5.200000000000000000e+01,5.600000000000000000e+01,5.200000000000000000e+01,5.000000000000000000e+01,4.600000000000000000e+01,3.700000000000000000e+01,2.600000000000000000e+01,3.000000000000000000e+01,3.100000000000000000e+01,3.600000000000000000e+01,3.900000000000000000e+01,5.100000000000000000e+01,5.300000000000000000e+01,4.300000000000000000e+01,5.800000000000000000e+01,1.220000000000000000e+02,1.400000000000000000e+02,1.120000000000000000e+02,1.380000000000000000e+02,1.710000000000000000e+02,1.810000000000000000e+02,1.710000000000000000e+02,1.480000000000000000e+02,1.460000000000000000e+02,1.300000000000000000e+02,1.220000000000000000e+02,1.380000000000000000e+02,1.340000000000000000e+02,1.430000000000000000e+02,1.360000000000000000e+02,1.210000000000000000e+02,1.160000000000000000e+02,1.130000000000000000e+02,1.390000000000000000e+02,1.630000000000000000e+02,1.700000000000000000e+02,1.750000000000000000e+02,1.860000000000000000e+02,1.820000000000000000e+02,1.830000000000000000e+02,2.120000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.120000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02),
(1.690000000000000000e+02,1.570000000000000000e+02,1.260000000000000000e+02,8.800000000000000000e+01,7.200000000000000000e+01,5.700000000000000000e+01,7.800000000000000000e+01,1.130000000000000000e+02,1.600000000000000000e+02,1.560000000000000000e+02,1.430000000000000000e+02,1.060000000000000000e+02,7.100000000000000000e+01,3.400000000000000000e+01,2.100000000000000000e+01,2.500000000000000000e+01,3.300000000000000000e+01,2.600000000000000000e+01,3.200000000000000000e+01,2.300000000000000000e+01,2.400000000000000000e+01,1.280000000000000000e+02,8.300000000000000000e+01,1.050000000000000000e+02,1.190000000000000000e+02,1.000000000000000000e+02,1.040000000000000000e+02,1.230000000000000000e+02,1.470000000000000000e+02,1.600000000000000000e+02,1.840000000000000000e+02,1.850000000000000000e+02,1.870000000000000000e+02,1.920000000000000000e+02,1.950000000000000000e+02,1.890000000000000000e+02,1.900000000000000000e+02,1.870000000000000000e+02,1.780000000000000000e+02,1.880000000000000000e+02,1.810000000000000000e+02,1.750000000000000000e+02,1.570000000000000000e+02,1.390000000000000000e+02,1.350000000000000000e+02,1.360000000000000000e+02,1.140000000000000000e+02,1.270000000000000000e+02,1.000000000000000000e+02,2.700000000000000000e+01,3.000000000000000000e+01,2.400000000000000000e+01,2.300000000000000000e+01,2.600000000000000000e+01,3.100000000000000000e+01,3.500000000000000000e+01,4.000000000000000000e+01,4.300000000000000000e+01,5.200000000000000000e+01,4.500000000000000000e+01,4.800000000000000000e+01,4.000000000000000000e+01,3.100000000000000000e+01,2.400000000000000000e+01,2.300000000000000000e+01,2.600000000000000000e+01,2.900000000000000000e+01,3.900000000000000000e+01,3.600000000000000000e+01,4.400000000000000000e+01,4.500000000000000000e+01,3.700000000000000000e+01,3.700000000000000000e+01,3.700000000000000000e+01,2.800000000000000000e+01,3.400000000000000000e+01,3.900000000000000000e+01,4.100000000000000000e+01,5.000000000000000000e+01,6.000000000000000000e+01,6.300000000000000000e+01,6.500000000000000000e+01,6.300000000000000000e+01,5.400000000000000000e+01,4.200000000000000000e+01,3.600000000000000000e+01,4.000000000000000000e+01,4.000000000000000000e+01,4.000000000000000000e+01,5.000000000000000000e+01,4.700000000000000000e+01,5.400000000000000000e+01,7.900000000000000000e+01,1.220000000000000000e+02,1.390000000000000000e+02,1.200000000000000000e+02,1.470000000000000000e+02,1.780000000000000000e+02,1.770000000000000000e+02,1.500000000000000000e+02,1.320000000000000000e+02,1.210000000000000000e+02,1.150000000000000000e+02,1.090000000000000000e+02,1.240000000000000000e+02,1.240000000000000000e+02,1.300000000000000000e+02,1.350000000000000000e+02,1.410000000000000000e+02,1.390000000000000000e+02,1.160000000000000000e+02,1.230000000000000000e+02,1.500000000000000000e+02,1.680000000000000000e+02,1.660000000000000000e+02,1.700000000000000000e+02,1.780000000000000000e+02,1.840000000000000000e+02,1.830000000000000000e+02,2.110000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02),
(1.680000000000000000e+02,1.550000000000000000e+02,1.310000000000000000e+02,9.200000000000000000e+01,7.000000000000000000e+01,5.300000000000000000e+01,7.700000000000000000e+01,1.120000000000000000e+02,1.540000000000000000e+02,1.530000000000000000e+02,1.350000000000000000e+02,1.050000000000000000e+02,6.700000000000000000e+01,3.600000000000000000e+01,2.400000000000000000e+01,2.800000000000000000e+01,2.700000000000000000e+01,2.600000000000000000e+01,2.900000000000000000e+01,2.900000000000000000e+01,2.900000000000000000e+01,1.250000000000000000e+02,1.010000000000000000e+02,1.220000000000000000e+02,1.140000000000000000e+02,9.300000000000000000e+01,1.100000000000000000e+02,1.400000000000000000e+02,1.490000000000000000e+02,1.780000000000000000e+02,1.820000000000000000e+02,1.810000000000000000e+02,1.850000000000000000e+02,1.890000000000000000e+02,1.940000000000000000e+02,1.790000000000000000e+02,1.780000000000000000e+02,1.810000000000000000e+02,1.730000000000000000e+02,1.900000000000000000e+02,1.740000000000000000e+02,1.710000000000000000e+02,1.740000000000000000e+02,1.530000000000000000e+02,1.310000000000000000e+02,1.250000000000000000e+02,1.300000000000000000e+02,1.160000000000000000e+02,1.320000000000000000e+02,4.900000000000000000e+01,5.300000000000000000e+01,6.200000000000000000e+01,4.600000000000000000e+01,5.800000000000000000e+01,6.400000000000000000e+01,6.600000000000000000e+01,7.400000000000000000e+01,6.500000000000000000e+01,8.100000000000000000e+01,7.200000000000000000e+01,8.200000000000000000e+01,7.300000000000000000e+01,7.400000000000000000e+01,6.700000000000000000e+01,6.400000000000000000e+01,6.700000000000000000e+01,6.900000000000000000e+01,7.000000000000000000e+01,7.800000000000000000e+01,7.800000000000000000e+01,7.700000000000000000e+01,7.900000000000000000e+01,8.500000000000000000e+01,8.000000000000000000e+01,7.800000000000000000e+01,8.400000000000000000e+01,8.600000000000000000e+01,9.000000000000000000e+01,9.300000000000000000e+01,9.700000000000000000e+01,1.040000000000000000e+02,1.100000000000000000e+02,1.040000000000000000e+02,9.800000000000000000e+01,9.600000000000000000e+01,9.100000000000000000e+01,9.400000000000000000e+01,9.100000000000000000e+01,8.900000000000000000e+01,9.300000000000000000e+01,7.600000000000000000e+01,1.110000000000000000e+02,1.310000000000000000e+02,1.490000000000000000e+02,1.450000000000000000e+02,1.580000000000000000e+02,1.810000000000000000e+02,1.670000000000000000e+02,1.610000000000000000e+02,1.530000000000000000e+02,1.410000000000000000e+02,1.410000000000000000e+02,1.210000000000000000e+02,1.150000000000000000e+02,1.260000000000000000e+02,1.460000000000000000e+02,1.440000000000000000e+02,1.450000000000000000e+02,1.460000000000000000e+02,1.340000000000000000e+02,1.300000000000000000e+02,1.390000000000000000e+02,1.660000000000000000e+02,1.720000000000000000e+02,1.750000000000000000e+02,1.760000000000000000e+02,1.840000000000000000e+02,1.870000000000000000e+02,1.860000000000000000e+02,2.110000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02),
(1.660000000000000000e+02,1.530000000000000000e+02,1.330000000000000000e+02,9.100000000000000000e+01,6.500000000000000000e+01,4.600000000000000000e+01,7.300000000000000000e+01,1.090000000000000000e+02,1.480000000000000000e+02,1.500000000000000000e+02,1.370000000000000000e+02,1.060000000000000000e+02,7.700000000000000000e+01,4.900000000000000000e+01,3.300000000000000000e+01,4.300000000000000000e+01,4.800000000000000000e+01,4.800000000000000000e+01,5.500000000000000000e+01,6.100000000000000000e+01,5.700000000000000000e+01,1.230000000000000000e+02,1.220000000000000000e+02,1.300000000000000000e+02,1.140000000000000000e+02,9.300000000000000000e+01,1.190000000000000000e+02,1.450000000000000000e+02,1.630000000000000000e+02,1.740000000000000000e+02,1.720000000000000000e+02,1.870000000000000000e+02,1.770000000000000000e+02,1.970000000000000000e+02,1.930000000000000000e+02,1.840000000000000000e+02,1.800000000000000000e+02,1.830000000000000000e+02,1.850000000000000000e+02,1.710000000000000000e+02,1.660000000000000000e+02,1.540000000000000000e+02,1.640000000000000000e+02,1.400000000000000000e+02,1.460000000000000000e+02,1.020000000000000000e+02,1.450000000000000000e+02,1.120000000000000000e+02,1.350000000000000000e+02,1.030000000000000000e+02,9.600000000000000000e+01,1.020000000000000000e+02,1.100000000000000000e+02,1.130000000000000000e+02,1.130000000000000000e+02,1.160000000000000000e+02,1.210000000000000000e+02,1.210000000000000000e+02,1.420000000000000000e+02,1.230000000000000000e+02,1.240000000000000000e+02,1.250000000000000000e+02,1.250000000000000000e+02,1.290000000000000000e+02,1.260000000000000000e+02,1.320000000000000000e+02,1.250000000000000000e+02,1.120000000000000000e+02,1.240000000000000000e+02,1.290000000000000000e+02,1.280000000000000000e+02,1.330000000000000000e+02,1.430000000000000000e+02,1.350000000000000000e+02,1.380000000000000000e+02,1.420000000000000000e+02,1.360000000000000000e+02,1.380000000000000000e+02,1.470000000000000000e+02,1.470000000000000000e+02,1.490000000000000000e+02,1.510000000000000000e+02,1.520000000000000000e+02,1.520000000000000000e+02,1.520000000000000000e+02,1.530000000000000000e+02,1.410000000000000000e+02,1.410000000000000000e+02,1.350000000000000000e+02,1.130000000000000000e+02,1.000000000000000000e+02,1.460000000000000000e+02,1.390000000000000000e+02,1.360000000000000000e+02,1.670000000000000000e+02,1.820000000000000000e+02,1.710000000000000000e+02,1.600000000000000000e+02,1.660000000000000000e+02,1.710000000000000000e+02,1.790000000000000000e+02,1.810000000000000000e+02,1.690000000000000000e+02,1.670000000000000000e+02,1.580000000000000000e+02,1.540000000000000000e+02,1.570000000000000000e+02,1.630000000000000000e+02,1.500000000000000000e+02,1.490000000000000000e+02,1.420000000000000000e+02,1.540000000000000000e+02,1.790000000000000000e+02,1.820000000000000000e+02,1.750000000000000000e+02,1.840000000000000000e+02,1.850000000000000000e+02,1.880000000000000000e+02,1.880000000000000000e+02,2.120000000000000000e+02,2.130000000000000000e+02,2.140000000000000000e+02,2.150000000000000000e+02,2.150000000000000000e+02,2.150000000000000000e+02,2.150000000000000000e+02,2.140000000000000000e+02,2.140000000000000000e+02),
(1.660000000000000000e+02,1.550000000000000000e+02,1.240000000000000000e+02,9.300000000000000000e+01,6.700000000000000000e+01,4.500000000000000000e+01,7.700000000000000000e+01,1.080000000000000000e+02,1.430000000000000000e+02,1.450000000000000000e+02,1.400000000000000000e+02,1.180000000000000000e+02,9.200000000000000000e+01,7.000000000000000000e+01,6.400000000000000000e+01,7.100000000000000000e+01,7.600000000000000000e+01,8.800000000000000000e+01,8.700000000000000000e+01,9.000000000000000000e+01,9.400000000000000000e+01,1.140000000000000000e+02,1.340000000000000000e+02,1.440000000000000000e+02,1.140000000000000000e+02,9.300000000000000000e+01,1.350000000000000000e+02,1.460000000000000000e+02,1.430000000000000000e+02,1.570000000000000000e+02,1.800000000000000000e+02,1.590000000000000000e+02,1.580000000000000000e+02,1.520000000000000000e+02,1.570000000000000000e+02,1.940000000000000000e+02,1.980000000000000000e+02,1.890000000000000000e+02,1.910000000000000000e+02,2.000000000000000000e+02,1.880000000000000000e+02,1.740000000000000000e+02,1.550000000000000000e+02,1.430000000000000000e+02,1.440000000000000000e+02,1.420000000000000000e+02,1.370000000000000000e+02,1.130000000000000000e+02,1.180000000000000000e+02,1.470000000000000000e+02,1.200000000000000000e+02,1.450000000000000000e+02,1.540000000000000000e+02,1.630000000000000000e+02,1.610000000000000000e+02,1.620000000000000000e+02,1.640000000000000000e+02,1.670000000000000000e+02,1.700000000000000000e+02,1.620000000000000000e+02,1.620000000000000000e+02,1.670000000000000000e+02,1.700000000000000000e+02,1.690000000000000000e+02,1.690000000000000000e+02,1.630000000000000000e+02,1.680000000000000000e+02,1.690000000000000000e+02,1.670000000000000000e+02,1.680000000000000000e+02,1.700000000000000000e+02,1.730000000000000000e+02,1.700000000000000000e+02,1.780000000000000000e+02,1.800000000000000000e+02,1.790000000000000000e+02,1.790000000000000000e+02,1.740000000000000000e+02,1.810000000000000000e+02,1.830000000000000000e+02,1.800000000000000000e+02,1.810000000000000000e+02,1.770000000000000000e+02,1.800000000000000000e+02,1.820000000000000000e+02,1.790000000000000000e+02,1.750000000000000000e+02,1.680000000000000000e+02,1.580000000000000000e+02,1.200000000000000000e+02,1.320000000000000000e+02,1.310000000000000000e+02,1.320000000000000000e+02,1.520000000000000000e+02,1.720000000000000000e+02,1.630000000000000000e+02,1.690000000000000000e+02,1.890000000000000000e+02,1.900000000000000000e+02,1.850000000000000000e+02,1.750000000000000000e+02,1.820000000000000000e+02,1.770000000000000000e+02,1.710000000000000000e+02,1.620000000000000000e+02,1.600000000000000000e+02,1.600000000000000000e+02,1.690000000000000000e+02,1.620000000000000000e+02,1.340000000000000000e+02,1.290000000000000000e+02,1.670000000000000000e+02,1.870000000000000000e+02,1.830000000000000000e+02,1.860000000000000000e+02,1.870000000000000000e+02,1.890000000000000000e+02,1.900000000000000000e+02,1.880000000000000000e+02,2.030000000000000000e+02,2.120000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.120000000000000000e+02,2.120000000000000000e+02),
(1.650000000000000000e+02,1.550000000000000000e+02,1.210000000000000000e+02,8.700000000000000000e+01,6.400000000000000000e+01,4.600000000000000000e+01,7.100000000000000000e+01,1.010000000000000000e+02,1.430000000000000000e+02,1.430000000000000000e+02,1.410000000000000000e+02,1.280000000000000000e+02,1.050000000000000000e+02,9.700000000000000000e+01,9.500000000000000000e+01,1.000000000000000000e+02,1.090000000000000000e+02,1.190000000000000000e+02,1.160000000000000000e+02,1.160000000000000000e+02,1.210000000000000000e+02,1.100000000000000000e+02,1.450000000000000000e+02,1.450000000000000000e+02,1.100000000000000000e+02,1.020000000000000000e+02,1.160000000000000000e+02,1.260000000000000000e+02,1.320000000000000000e+02,1.620000000000000000e+02,1.470000000000000000e+02,1.660000000000000000e+02,1.810000000000000000e+02,1.810000000000000000e+02,1.800000000000000000e+02,1.660000000000000000e+02,1.790000000000000000e+02,1.970000000000000000e+02,1.880000000000000000e+02,1.840000000000000000e+02,1.870000000000000000e+02,1.780000000000000000e+02,1.580000000000000000e+02,1.380000000000000000e+02,1.470000000000000000e+02,1.190000000000000000e+02,1.240000000000000000e+02,9.100000000000000000e+01,1.080000000000000000e+02,1.270000000000000000e+02,1.490000000000000000e+02,1.670000000000000000e+02,1.860000000000000000e+02,1.840000000000000000e+02,1.880000000000000000e+02,1.870000000000000000e+02,1.870000000000000000e+02,1.880000000000000000e+02,1.970000000000000000e+02,1.900000000000000000e+02,1.910000000000000000e+02,1.930000000000000000e+02,1.900000000000000000e+02,1.890000000000000000e+02,1.930000000000000000e+02,1.900000000000000000e+02,1.870000000000000000e+02,1.950000000000000000e+02,1.910000000000000000e+02,1.910000000000000000e+02,1.920000000000000000e+02,1.920000000000000000e+02,1.970000000000000000e+02,1.950000000000000000e+02,1.950000000000000000e+02,1.960000000000000000e+02,1.960000000000000000e+02,1.940000000000000000e+02,1.990000000000000000e+02,1.980000000000000000e+02,1.970000000000000000e+02,1.990000000000000000e+02,1.990000000000000000e+02,1.990000000000000000e+02,1.970000000000000000e+02,1.950000000000000000e+02,1.940000000000000000e+02,1.800000000000000000e+02,1.580000000000000000e+02,1.380000000000000000e+02,1.490000000000000000e+02,1.630000000000000000e+02,1.510000000000000000e+02,1.820000000000000000e+02,1.840000000000000000e+02,1.830000000000000000e+02,1.790000000000000000e+02,1.770000000000000000e+02,1.610000000000000000e+02,1.550000000000000000e+02,1.500000000000000000e+02,1.530000000000000000e+02,1.550000000000000000e+02,1.660000000000000000e+02,1.690000000000000000e+02,1.700000000000000000e+02,1.650000000000000000e+02,1.630000000000000000e+02,1.500000000000000000e+02,1.350000000000000000e+02,1.540000000000000000e+02,1.830000000000000000e+02,1.910000000000000000e+02,1.910000000000000000e+02,1.920000000000000000e+02,1.900000000000000000e+02,1.890000000000000000e+02,1.920000000000000000e+02,1.920000000000000000e+02,1.920000000000000000e+02,1.970000000000000000e+02,2.080000000000000000e+02,2.100000000000000000e+02,2.100000000000000000e+02,2.100000000000000000e+02,2.090000000000000000e+02,2.090000000000000000e+02,2.070000000000000000e+02),
(1.640000000000000000e+02,1.540000000000000000e+02,1.270000000000000000e+02,9.400000000000000000e+01,6.600000000000000000e+01,4.700000000000000000e+01,6.900000000000000000e+01,9.900000000000000000e+01,1.420000000000000000e+02,1.470000000000000000e+02,1.470000000000000000e+02,1.390000000000000000e+02,1.270000000000000000e+02,1.110000000000000000e+02,1.210000000000000000e+02,1.330000000000000000e+02,1.330000000000000000e+02,1.430000000000000000e+02,1.450000000000000000e+02,1.430000000000000000e+02,1.470000000000000000e+02,1.200000000000000000e+02,1.450000000000000000e+02,1.570000000000000000e+02,1.220000000000000000e+02,9.800000000000000000e+01,1.150000000000000000e+02,1.220000000000000000e+02,1.100000000000000000e+02,1.310000000000000000e+02,1.250000000000000000e+02,1.290000000000000000e+02,1.380000000000000000e+02,1.490000000000000000e+02,1.800000000000000000e+02,1.510000000000000000e+02,1.580000000000000000e+02,1.710000000000000000e+02,1.740000000000000000e+02,1.950000000000000000e+02,1.800000000000000000e+02,1.690000000000000000e+02,1.550000000000000000e+02,1.540000000000000000e+02,1.380000000000000000e+02,1.360000000000000000e+02,1.140000000000000000e+02,8.600000000000000000e+01,8.600000000000000000e+01,9.000000000000000000e+01,1.560000000000000000e+02,1.550000000000000000e+02,1.960000000000000000e+02,1.970000000000000000e+02,1.970000000000000000e+02,2.020000000000000000e+02,2.000000000000000000e+02,2.020000000000000000e+02,2.010000000000000000e+02,2.010000000000000000e+02,2.030000000000000000e+02,2.020000000000000000e+02,2.040000000000000000e+02,2.050000000000000000e+02,2.030000000000000000e+02,2.030000000000000000e+02,1.970000000000000000e+02,2.020000000000000000e+02,2.030000000000000000e+02,2.030000000000000000e+02,2.040000000000000000e+02,2.040000000000000000e+02,2.040000000000000000e+02,2.050000000000000000e+02,2.020000000000000000e+02,2.030000000000000000e+02,2.040000000000000000e+02,2.060000000000000000e+02,2.050000000000000000e+02,2.030000000000000000e+02,2.020000000000000000e+02,2.030000000000000000e+02,2.050000000000000000e+02,2.050000000000000000e+02,2.020000000000000000e+02,1.980000000000000000e+02,1.970000000000000000e+02,1.620000000000000000e+02,1.530000000000000000e+02,1.470000000000000000e+02,1.690000000000000000e+02,1.570000000000000000e+02,1.640000000000000000e+02,1.750000000000000000e+02,1.650000000000000000e+02,1.640000000000000000e+02,1.530000000000000000e+02,1.590000000000000000e+02,1.720000000000000000e+02,1.670000000000000000e+02,1.720000000000000000e+02,1.750000000000000000e+02,1.740000000000000000e+02,1.670000000000000000e+02,1.700000000000000000e+02,1.780000000000000000e+02,1.800000000000000000e+02,1.680000000000000000e+02,1.530000000000000000e+02,1.420000000000000000e+02,1.650000000000000000e+02,1.930000000000000000e+02,1.930000000000000000e+02,1.930000000000000000e+02,1.960000000000000000e+02,1.950000000000000000e+02,1.950000000000000000e+02,1.920000000000000000e+02,1.940000000000000000e+02,1.910000000000000000e+02,1.910000000000000000e+02,1.900000000000000000e+02,1.910000000000000000e+02,1.910000000000000000e+02,1.910000000000000000e+02,1.900000000000000000e+02,1.910000000000000000e+02,1.900000000000000000e+02),
(1.610000000000000000e+02,1.510000000000000000e+02,1.310000000000000000e+02,8.500000000000000000e+01,6.300000000000000000e+01,4.200000000000000000e+01,6.700000000000000000e+01,9.700000000000000000e+01,1.370000000000000000e+02,1.500000000000000000e+02,1.490000000000000000e+02,1.480000000000000000e+02,1.410000000000000000e+02,1.330000000000000000e+02,1.430000000000000000e+02,1.500000000000000000e+02,1.530000000000000000e+02,1.590000000000000000e+02,1.600000000000000000e+02,1.640000000000000000e+02,1.630000000000000000e+02,1.210000000000000000e+02,1.550000000000000000e+02,1.620000000000000000e+02,1.230000000000000000e+02,1.080000000000000000e+02,1.210000000000000000e+02,1.180000000000000000e+02,1.140000000000000000e+02,1.180000000000000000e+02,1.160000000000000000e+02,1.160000000000000000e+02,1.220000000000000000e+02,1.330000000000000000e+02,1.580000000000000000e+02,1.620000000000000000e+02,1.530000000000000000e+02,1.510000000000000000e+02,1.550000000000000000e+02,1.700000000000000000e+02,1.840000000000000000e+02,1.890000000000000000e+02,1.630000000000000000e+02,1.430000000000000000e+02,1.190000000000000000e+02,1.140000000000000000e+02,6.300000000000000000e+01,8.400000000000000000e+01,8.500000000000000000e+01,8.100000000000000000e+01,1.190000000000000000e+02,1.640000000000000000e+02,1.720000000000000000e+02,1.920000000000000000e+02,1.990000000000000000e+02,2.050000000000000000e+02,2.030000000000000000e+02,2.030000000000000000e+02,2.030000000000000000e+02,2.050000000000000000e+02,2.050000000000000000e+02,2.040000000000000000e+02,2.050000000000000000e+02,2.050000000000000000e+02,2.060000000000000000e+02,2.050000000000000000e+02,2.030000000000000000e+02,2.030000000000000000e+02,2.040000000000000000e+02,2.040000000000000000e+02,2.050000000000000000e+02,2.050000000000000000e+02,2.060000000000000000e+02,2.050000000000000000e+02,2.040000000000000000e+02,2.040000000000000000e+02,2.050000000000000000e+02,2.050000000000000000e+02,2.040000000000000000e+02,2.030000000000000000e+02,2.030000000000000000e+02,2.030000000000000000e+02,2.030000000000000000e+02,2.030000000000000000e+02,2.010000000000000000e+02,1.930000000000000000e+02,1.720000000000000000e+02,1.510000000000000000e+02,1.520000000000000000e+02,1.440000000000000000e+02,1.520000000000000000e+02,1.580000000000000000e+02,1.810000000000000000e+02,1.880000000000000000e+02,1.890000000000000000e+02,1.860000000000000000e+02,1.920000000000000000e+02,1.960000000000000000e+02,1.980000000000000000e+02,1.930000000000000000e+02,1.890000000000000000e+02,1.830000000000000000e+02,1.670000000000000000e+02,1.690000000000000000e+02,1.760000000000000000e+02,1.790000000000000000e+02,1.770000000000000000e+02,1.700000000000000000e+02,1.480000000000000000e+02,1.370000000000000000e+02,1.790000000000000000e+02,1.900000000000000000e+02,1.920000000000000000e+02,1.920000000000000000e+02,1.890000000000000000e+02,1.880000000000000000e+02,1.870000000000000000e+02,1.870000000000000000e+02,1.850000000000000000e+02,1.870000000000000000e+02,1.850000000000000000e+02,1.850000000000000000e+02,1.840000000000000000e+02,1.850000000000000000e+02,1.860000000000000000e+02,1.810000000000000000e+02,1.830000000000000000e+02,1.810000000000000000e+02),
(1.580000000000000000e+02,1.510000000000000000e+02,1.190000000000000000e+02,8.600000000000000000e+01,6.100000000000000000e+01,4.100000000000000000e+01,6.800000000000000000e+01,9.600000000000000000e+01,1.400000000000000000e+02,1.440000000000000000e+02,1.470000000000000000e+02,1.440000000000000000e+02,1.440000000000000000e+02,1.390000000000000000e+02,1.460000000000000000e+02,1.510000000000000000e+02,1.530000000000000000e+02,1.550000000000000000e+02,1.600000000000000000e+02,1.660000000000000000e+02,1.690000000000000000e+02,1.430000000000000000e+02,1.400000000000000000e+02,1.590000000000000000e+02,1.360000000000000000e+02,1.080000000000000000e+02,1.170000000000000000e+02,1.190000000000000000e+02,1.250000000000000000e+02,1.300000000000000000e+02,1.320000000000000000e+02,1.240000000000000000e+02,1.400000000000000000e+02,1.230000000000000000e+02,1.190000000000000000e+02,1.240000000000000000e+02,1.250000000000000000e+02,1.240000000000000000e+02,1.130000000000000000e+02,1.460000000000000000e+02,1.550000000000000000e+02,1.800000000000000000e+02,1.770000000000000000e+02,1.400000000000000000e+02,1.230000000000000000e+02,1.160000000000000000e+02,8.100000000000000000e+01,7.600000000000000000e+01,5.900000000000000000e+01,5.700000000000000000e+01,7.400000000000000000e+01,1.280000000000000000e+02,1.680000000000000000e+02,1.580000000000000000e+02,1.880000000000000000e+02,1.920000000000000000e+02,1.980000000000000000e+02,2.010000000000000000e+02,2.000000000000000000e+02,2.010000000000000000e+02,2.010000000000000000e+02,2.020000000000000000e+02,2.030000000000000000e+02,2.030000000000000000e+02,2.010000000000000000e+02,2.040000000000000000e+02,2.000000000000000000e+02,2.030000000000000000e+02,2.030000000000000000e+02,2.030000000000000000e+02,2.030000000000000000e+02,2.030000000000000000e+02,2.030000000000000000e+02,2.020000000000000000e+02,2.040000000000000000e+02,2.040000000000000000e+02,2.030000000000000000e+02,2.030000000000000000e+02,2.010000000000000000e+02,2.000000000000000000e+02,1.990000000000000000e+02,1.990000000000000000e+02,1.990000000000000000e+02,1.960000000000000000e+02,1.870000000000000000e+02,1.620000000000000000e+02,1.690000000000000000e+02,1.310000000000000000e+02,1.440000000000000000e+02,1.580000000000000000e+02,1.600000000000000000e+02,1.740000000000000000e+02,1.750000000000000000e+02,1.850000000000000000e+02,1.900000000000000000e+02,1.890000000000000000e+02,1.980000000000000000e+02,1.990000000000000000e+02,1.980000000000000000e+02,1.990000000000000000e+02,2.020000000000000000e+02,1.960000000000000000e+02,1.890000000000000000e+02,1.910000000000000000e+02,1.890000000000000000e+02,1.920000000000000000e+02,1.830000000000000000e+02,1.670000000000000000e+02,1.480000000000000000e+02,1.490000000000000000e+02,1.780000000000000000e+02,1.840000000000000000e+02,1.850000000000000000e+02,1.850000000000000000e+02,1.830000000000000000e+02,1.850000000000000000e+02,1.810000000000000000e+02,1.810000000000000000e+02,1.830000000000000000e+02,1.810000000000000000e+02,1.820000000000000000e+02,1.820000000000000000e+02,1.820000000000000000e+02,1.750000000000000000e+02,1.730000000000000000e+02,1.720000000000000000e+02,1.740000000000000000e+02,1.730000000000000000e+02),
(1.600000000000000000e+02,1.420000000000000000e+02,1.180000000000000000e+02,8.100000000000000000e+01,5.900000000000000000e+01,4.000000000000000000e+01,6.900000000000000000e+01,9.500000000000000000e+01,1.350000000000000000e+02,1.430000000000000000e+02,1.450000000000000000e+02,1.480000000000000000e+02,1.430000000000000000e+02,1.350000000000000000e+02,1.370000000000000000e+02,1.460000000000000000e+02,1.510000000000000000e+02,1.570000000000000000e+02,1.600000000000000000e+02,1.610000000000000000e+02,1.610000000000000000e+02,1.310000000000000000e+02,1.460000000000000000e+02,1.530000000000000000e+02,1.560000000000000000e+02,1.070000000000000000e+02,1.060000000000000000e+02,1.220000000000000000e+02,1.170000000000000000e+02,1.160000000000000000e+02,1.170000000000000000e+02,1.180000000000000000e+02,1.110000000000000000e+02,1.160000000000000000e+02,1.240000000000000000e+02,1.210000000000000000e+02,1.190000000000000000e+02,1.310000000000000000e+02,1.370000000000000000e+02,1.560000000000000000e+02,1.630000000000000000e+02,1.660000000000000000e+02,1.690000000000000000e+02,1.620000000000000000e+02,1.380000000000000000e+02,1.150000000000000000e+02,8.700000000000000000e+01,6.800000000000000000e+01,6.600000000000000000e+01,7.800000000000000000e+01,8.700000000000000000e+01,1.260000000000000000e+02,1.750000000000000000e+02,1.730000000000000000e+02,1.490000000000000000e+02,1.580000000000000000e+02,1.890000000000000000e+02,1.950000000000000000e+02,1.940000000000000000e+02,1.970000000000000000e+02,1.930000000000000000e+02,1.990000000000000000e+02,1.970000000000000000e+02,2.020000000000000000e+02,1.990000000000000000e+02,2.010000000000000000e+02,2.040000000000000000e+02,2.020000000000000000e+02,2.020000000000000000e+02,1.990000000000000000e+02,1.990000000000000000e+02,2.050000000000000000e+02,2.020000000000000000e+02,1.980000000000000000e+02,2.010000000000000000e+02,2.020000000000000000e+02,1.980000000000000000e+02,1.980000000000000000e+02,1.960000000000000000e+02,1.950000000000000000e+02,1.950000000000000000e+02,1.930000000000000000e+02,1.880000000000000000e+02,1.690000000000000000e+02,1.370000000000000000e+02,1.610000000000000000e+02,1.470000000000000000e+02,1.470000000000000000e+02,1.370000000000000000e+02,1.490000000000000000e+02,1.630000000000000000e+02,1.840000000000000000e+02,1.990000000000000000e+02,2.050000000000000000e+02,1.930000000000000000e+02,2.010000000000000000e+02,1.990000000000000000e+02,1.970000000000000000e+02,1.980000000000000000e+02,1.950000000000000000e+02,1.930000000000000000e+02,1.930000000000000000e+02,1.980000000000000000e+02,2.010000000000000000e+02,2.000000000000000000e+02,1.950000000000000000e+02,1.860000000000000000e+02,1.620000000000000000e+02,1.370000000000000000e+02,1.530000000000000000e+02,1.740000000000000000e+02,1.750000000000000000e+02,1.750000000000000000e+02,1.730000000000000000e+02,1.760000000000000000e+02,1.750000000000000000e+02,1.770000000000000000e+02,1.710000000000000000e+02,1.700000000000000000e+02,1.750000000000000000e+02,1.680000000000000000e+02,1.660000000000000000e+02,1.660000000000000000e+02,1.660000000000000000e+02,1.610000000000000000e+02,1.610000000000000000e+02,1.550000000000000000e+02,1.520000000000000000e+02),
(1.550000000000000000e+02,1.410000000000000000e+02,1.160000000000000000e+02,7.800000000000000000e+01,5.200000000000000000e+01,3.500000000000000000e+01,6.900000000000000000e+01,9.200000000000000000e+01,1.360000000000000000e+02,1.450000000000000000e+02,1.410000000000000000e+02,1.460000000000000000e+02,1.370000000000000000e+02,1.380000000000000000e+02,1.370000000000000000e+02,1.360000000000000000e+02,1.470000000000000000e+02,1.550000000000000000e+02,1.530000000000000000e+02,1.620000000000000000e+02,1.440000000000000000e+02,1.600000000000000000e+02,1.470000000000000000e+02,1.510000000000000000e+02,1.650000000000000000e+02,1.340000000000000000e+02,1.220000000000000000e+02,1.360000000000000000e+02,1.370000000000000000e+02,1.430000000000000000e+02,1.400000000000000000e+02,1.300000000000000000e+02,1.280000000000000000e+02,1.200000000000000000e+02,1.130000000000000000e+02,1.170000000000000000e+02,1.130000000000000000e+02,1.330000000000000000e+02,1.590000000000000000e+02,1.640000000000000000e+02,1.660000000000000000e+02,1.680000000000000000e+02,1.730000000000000000e+02,1.310000000000000000e+02,1.030000000000000000e+02,9.400000000000000000e+01,8.900000000000000000e+01,5.600000000000000000e+01,7.300000000000000000e+01,9.800000000000000000e+01,8.800000000000000000e+01,1.120000000000000000e+02,1.580000000000000000e+02,1.850000000000000000e+02,1.760000000000000000e+02,8.300000000000000000e+01,1.510000000000000000e+02,1.500000000000000000e+02,1.810000000000000000e+02,1.850000000000000000e+02,1.620000000000000000e+02,1.830000000000000000e+02,1.830000000000000000e+02,1.900000000000000000e+02,1.940000000000000000e+02,1.820000000000000000e+02,1.920000000000000000e+02,1.910000000000000000e+02,1.890000000000000000e+02,1.890000000000000000e+02,1.930000000000000000e+02,1.870000000000000000e+02,1.870000000000000000e+02,1.880000000000000000e+02,1.870000000000000000e+02,1.830000000000000000e+02,1.770000000000000000e+02,1.800000000000000000e+02,1.790000000000000000e+02,1.740000000000000000e+02,1.690000000000000000e+02,1.480000000000000000e+02,1.140000000000000000e+02,6.900000000000000000e+01,1.320000000000000000e+02,1.230000000000000000e+02,1.200000000000000000e+02,1.150000000000000000e+02,1.370000000000000000e+02,1.490000000000000000e+02,1.820000000000000000e+02,1.950000000000000000e+02,2.000000000000000000e+02,2.010000000000000000e+02,1.910000000000000000e+02,1.920000000000000000e+02,1.970000000000000000e+02,1.990000000000000000e+02,1.980000000000000000e+02,1.980000000000000000e+02,1.990000000000000000e+02,1.920000000000000000e+02,1.930000000000000000e+02,1.970000000000000000e+02,1.990000000000000000e+02,1.940000000000000000e+02,1.860000000000000000e+02,1.540000000000000000e+02,1.370000000000000000e+02,1.440000000000000000e+02,1.490000000000000000e+02,1.510000000000000000e+02,1.470000000000000000e+02,1.460000000000000000e+02,1.460000000000000000e+02,1.440000000000000000e+02,1.370000000000000000e+02,1.390000000000000000e+02,1.380000000000000000e+02,1.420000000000000000e+02,1.340000000000000000e+02,1.360000000000000000e+02,1.370000000000000000e+02,1.310000000000000000e+02,1.270000000000000000e+02,1.240000000000000000e+02,1.200000000000000000e+02,1.140000000000000000e+02),
(1.500000000000000000e+02,1.380000000000000000e+02,1.090000000000000000e+02,7.500000000000000000e+01,5.000000000000000000e+01,3.400000000000000000e+01,6.100000000000000000e+01,9.100000000000000000e+01,1.320000000000000000e+02,1.410000000000000000e+02,1.470000000000000000e+02,1.380000000000000000e+02,1.300000000000000000e+02,1.150000000000000000e+02,1.160000000000000000e+02,1.290000000000000000e+02,1.310000000000000000e+02,1.280000000000000000e+02,1.310000000000000000e+02,1.400000000000000000e+02,9.900000000000000000e+01,1.560000000000000000e+02,1.410000000000000000e+02,1.470000000000000000e+02,1.560000000000000000e+02,1.680000000000000000e+02,1.250000000000000000e+02,1.260000000000000000e+02,1.390000000000000000e+02,1.480000000000000000e+02,1.470000000000000000e+02,1.470000000000000000e+02,1.370000000000000000e+02,1.320000000000000000e+02,1.320000000000000000e+02,1.430000000000000000e+02,1.500000000000000000e+02,1.460000000000000000e+02,1.320000000000000000e+02,1.510000000000000000e+02,1.850000000000000000e+02,1.840000000000000000e+02,1.810000000000000000e+02,1.700000000000000000e+02,1.620000000000000000e+02,9.500000000000000000e+01,9.800000000000000000e+01,9.100000000000000000e+01,7.700000000000000000e+01,7.700000000000000000e+01,9.000000000000000000e+01,8.800000000000000000e+01,1.420000000000000000e+02,1.450000000000000000e+02,1.530000000000000000e+02,1.250000000000000000e+02,5.600000000000000000e+01,7.000000000000000000e+01,1.150000000000000000e+02,1.320000000000000000e+02,1.080000000000000000e+02,1.450000000000000000e+02,1.290000000000000000e+02,1.560000000000000000e+02,1.700000000000000000e+02,1.490000000000000000e+02,1.740000000000000000e+02,1.700000000000000000e+02,1.700000000000000000e+02,1.700000000000000000e+02,1.620000000000000000e+02,1.710000000000000000e+02,1.660000000000000000e+02,1.610000000000000000e+02,1.610000000000000000e+02,1.580000000000000000e+02,1.320000000000000000e+02,1.410000000000000000e+02,1.280000000000000000e+02,1.190000000000000000e+02,1.100000000000000000e+02,7.600000000000000000e+01,4.200000000000000000e+01,1.060000000000000000e+02,1.350000000000000000e+02,1.090000000000000000e+02,9.800000000000000000e+01,1.080000000000000000e+02,1.250000000000000000e+02,1.660000000000000000e+02,1.840000000000000000e+02,1.940000000000000000e+02,1.890000000000000000e+02,1.720000000000000000e+02,1.760000000000000000e+02,1.770000000000000000e+02,1.800000000000000000e+02,1.890000000000000000e+02,1.850000000000000000e+02,1.810000000000000000e+02,1.910000000000000000e+02,1.850000000000000000e+02,1.920000000000000000e+02,1.980000000000000000e+02,1.980000000000000000e+02,1.910000000000000000e+02,1.800000000000000000e+02,1.580000000000000000e+02,1.350000000000000000e+02,1.250000000000000000e+02,1.110000000000000000e+02,1.110000000000000000e+02,1.130000000000000000e+02,1.120000000000000000e+02,1.060000000000000000e+02,1.050000000000000000e+02,1.050000000000000000e+02,1.050000000000000000e+02,1.000000000000000000e+02,9.900000000000000000e+01,9.700000000000000000e+01,9.700000000000000000e+01,9.600000000000000000e+01,9.100000000000000000e+01,8.800000000000000000e+01,8.500000000000000000e+01,8.300000000000000000e+01,7.500000000000000000e+01),
(1.460000000000000000e+02,1.270000000000000000e+02,9.900000000000000000e+01,6.600000000000000000e+01,4.900000000000000000e+01,3.500000000000000000e+01,6.000000000000000000e+01,9.200000000000000000e+01,1.260000000000000000e+02,1.380000000000000000e+02,1.330000000000000000e+02,1.190000000000000000e+02,1.040000000000000000e+02,8.300000000000000000e+01,8.800000000000000000e+01,9.200000000000000000e+01,9.600000000000000000e+01,1.010000000000000000e+02,1.030000000000000000e+02,9.400000000000000000e+01,4.500000000000000000e+01,1.890000000000000000e+02,1.430000000000000000e+02,1.450000000000000000e+02,1.570000000000000000e+02,1.670000000000000000e+02,1.530000000000000000e+02,1.400000000000000000e+02,1.430000000000000000e+02,1.450000000000000000e+02,1.470000000000000000e+02,1.450000000000000000e+02,1.220000000000000000e+02,1.380000000000000000e+02,1.340000000000000000e+02,1.300000000000000000e+02,1.240000000000000000e+02,1.390000000000000000e+02,1.470000000000000000e+02,1.510000000000000000e+02,1.490000000000000000e+02,1.790000000000000000e+02,1.870000000000000000e+02,1.670000000000000000e+02,1.580000000000000000e+02,1.150000000000000000e+02,1.100000000000000000e+02,1.100000000000000000e+02,9.400000000000000000e+01,1.250000000000000000e+02,1.170000000000000000e+02,1.470000000000000000e+02,1.440000000000000000e+02,1.490000000000000000e+02,1.340000000000000000e+02,1.510000000000000000e+02,9.500000000000000000e+01,9.600000000000000000e+01,4.900000000000000000e+01,6.400000000000000000e+01,9.600000000000000000e+01,5.600000000000000000e+01,2.500000000000000000e+01,3.300000000000000000e+01,8.400000000000000000e+01,5.600000000000000000e+01,1.110000000000000000e+02,1.120000000000000000e+02,1.130000000000000000e+02,1.170000000000000000e+02,1.140000000000000000e+02,1.220000000000000000e+02,1.220000000000000000e+02,1.150000000000000000e+02,1.080000000000000000e+02,1.020000000000000000e+02,7.400000000000000000e+01,7.200000000000000000e+01,5.700000000000000000e+01,5.800000000000000000e+01,3.700000000000000000e+01,1.700000000000000000e+01,8.600000000000000000e+01,1.770000000000000000e+02,1.390000000000000000e+02,1.170000000000000000e+02,5.300000000000000000e+01,9.000000000000000000e+01,1.380000000000000000e+02,1.680000000000000000e+02,1.750000000000000000e+02,1.880000000000000000e+02,1.950000000000000000e+02,1.890000000000000000e+02,1.960000000000000000e+02,1.920000000000000000e+02,1.930000000000000000e+02,1.900000000000000000e+02,1.740000000000000000e+02,1.420000000000000000e+02,1.510000000000000000e+02,1.770000000000000000e+02,1.890000000000000000e+02,1.980000000000000000e+02,1.990000000000000000e+02,1.850000000000000000e+02,1.740000000000000000e+02,1.540000000000000000e+02,1.260000000000000000e+02,7.400000000000000000e+01,6.600000000000000000e+01,6.600000000000000000e+01,6.400000000000000000e+01,6.200000000000000000e+01,6.400000000000000000e+01,7.400000000000000000e+01,6.300000000000000000e+01,5.600000000000000000e+01,4.900000000000000000e+01,5.300000000000000000e+01,4.900000000000000000e+01,4.600000000000000000e+01,4.300000000000000000e+01,4.700000000000000000e+01,4.200000000000000000e+01,3.900000000000000000e+01,3.600000000000000000e+01,3.500000000000000000e+01),
(1.390000000000000000e+02,1.270000000000000000e+02,1.000000000000000000e+02,6.800000000000000000e+01,5.100000000000000000e+01,3.800000000000000000e+01,6.300000000000000000e+01,8.600000000000000000e+01,1.320000000000000000e+02,1.280000000000000000e+02,1.210000000000000000e+02,9.900000000000000000e+01,8.000000000000000000e+01,5.900000000000000000e+01,5.200000000000000000e+01,5.600000000000000000e+01,5.900000000000000000e+01,5.700000000000000000e+01,6.200000000000000000e+01,7.000000000000000000e+01,3.500000000000000000e+01,1.800000000000000000e+02,1.460000000000000000e+02,1.530000000000000000e+02,1.570000000000000000e+02,1.610000000000000000e+02,1.620000000000000000e+02,1.500000000000000000e+02,1.520000000000000000e+02,1.590000000000000000e+02,1.550000000000000000e+02,1.520000000000000000e+02,1.190000000000000000e+02,1.350000000000000000e+02,1.470000000000000000e+02,1.260000000000000000e+02,1.170000000000000000e+02,1.390000000000000000e+02,1.640000000000000000e+02,1.420000000000000000e+02,1.260000000000000000e+02,1.770000000000000000e+02,1.900000000000000000e+02,1.640000000000000000e+02,1.450000000000000000e+02,1.320000000000000000e+02,1.370000000000000000e+02,1.160000000000000000e+02,1.140000000000000000e+02,1.240000000000000000e+02,1.560000000000000000e+02,1.380000000000000000e+02,8.500000000000000000e+01,9.200000000000000000e+01,7.700000000000000000e+01,8.600000000000000000e+01,1.040000000000000000e+02,1.070000000000000000e+02,1.200000000000000000e+02,7.500000000000000000e+01,1.350000000000000000e+02,5.000000000000000000e+01,5.000000000000000000e+00,1.200000000000000000e+01,3.000000000000000000e+00,6.000000000000000000e+00,1.100000000000000000e+01,2.600000000000000000e+01,2.600000000000000000e+01,3.600000000000000000e+01,5.900000000000000000e+01,5.700000000000000000e+01,6.800000000000000000e+01,5.200000000000000000e+01,5.100000000000000000e+01,5.100000000000000000e+01,5.300000000000000000e+01,4.400000000000000000e+01,4.200000000000000000e+01,2.300000000000000000e+01,1.300000000000000000e+01,2.500000000000000000e+01,7.100000000000000000e+01,1.750000000000000000e+02,1.230000000000000000e+02,1.120000000000000000e+02,4.100000000000000000e+01,6.900000000000000000e+01,1.050000000000000000e+02,1.240000000000000000e+02,1.530000000000000000e+02,1.860000000000000000e+02,1.740000000000000000e+02,1.900000000000000000e+02,1.940000000000000000e+02,1.940000000000000000e+02,2.000000000000000000e+02,1.990000000000000000e+02,2.010000000000000000e+02,1.960000000000000000e+02,1.840000000000000000e+02,1.780000000000000000e+02,1.920000000000000000e+02,2.010000000000000000e+02,1.990000000000000000e+02,1.900000000000000000e+02,1.800000000000000000e+02,1.510000000000000000e+02,7.400000000000000000e+01,2.100000000000000000e+01,2.500000000000000000e+01,3.200000000000000000e+01,3.600000000000000000e+01,2.900000000000000000e+01,2.000000000000000000e+01,1.400000000000000000e+01,1.600000000000000000e+01,1.500000000000000000e+01,1.600000000000000000e+01,1.500000000000000000e+01,1.200000000000000000e+01,1.200000000000000000e+01,1.300000000000000000e+01,1.100000000000000000e+01,1.000000000000000000e+01,1.000000000000000000e+01,9.000000000000000000e+00,9.000000000000000000e+00),
(1.440000000000000000e+02,1.260000000000000000e+02,9.400000000000000000e+01,6.600000000000000000e+01,5.000000000000000000e+01,3.700000000000000000e+01,6.400000000000000000e+01,8.700000000000000000e+01,1.280000000000000000e+02,1.260000000000000000e+02,1.170000000000000000e+02,8.500000000000000000e+01,6.100000000000000000e+01,2.900000000000000000e+01,1.700000000000000000e+01,2.200000000000000000e+01,2.300000000000000000e+01,2.200000000000000000e+01,2.500000000000000000e+01,3.900000000000000000e+01,3.600000000000000000e+01,1.560000000000000000e+02,1.640000000000000000e+02,1.770000000000000000e+02,1.510000000000000000e+02,1.660000000000000000e+02,1.720000000000000000e+02,1.660000000000000000e+02,1.680000000000000000e+02,1.730000000000000000e+02,1.590000000000000000e+02,1.570000000000000000e+02,1.290000000000000000e+02,1.310000000000000000e+02,1.450000000000000000e+02,1.510000000000000000e+02,1.470000000000000000e+02,1.530000000000000000e+02,1.860000000000000000e+02,1.730000000000000000e+02,1.640000000000000000e+02,1.860000000000000000e+02,1.910000000000000000e+02,1.690000000000000000e+02,1.520000000000000000e+02,1.350000000000000000e+02,1.430000000000000000e+02,1.520000000000000000e+02,1.420000000000000000e+02,1.730000000000000000e+02,1.620000000000000000e+02,1.540000000000000000e+02,6.500000000000000000e+01,8.700000000000000000e+01,8.700000000000000000e+01,5.100000000000000000e+01,1.080000000000000000e+02,6.800000000000000000e+01,9.200000000000000000e+01,8.800000000000000000e+01,1.430000000000000000e+02,7.900000000000000000e+01,2.700000000000000000e+01,4.200000000000000000e+01,4.000000000000000000e+00,4.000000000000000000e+00,5.000000000000000000e+00,1.000000000000000000e+01,7.000000000000000000e+00,9.000000000000000000e+00,1.600000000000000000e+01,1.700000000000000000e+01,2.100000000000000000e+01,3.200000000000000000e+01,4.000000000000000000e+01,6.400000000000000000e+01,7.500000000000000000e+01,7.500000000000000000e+01,5.300000000000000000e+01,3.900000000000000000e+01,3.000000000000000000e+01,5.200000000000000000e+01,8.000000000000000000e+01,1.620000000000000000e+02,1.080000000000000000e+02,1.410000000000000000e+02,5.300000000000000000e+01,7.300000000000000000e+01,1.020000000000000000e+02,1.300000000000000000e+02,1.720000000000000000e+02,1.820000000000000000e+02,1.780000000000000000e+02,1.890000000000000000e+02,1.840000000000000000e+02,1.690000000000000000e+02,1.780000000000000000e+02,1.810000000000000000e+02,1.870000000000000000e+02,1.890000000000000000e+02,1.920000000000000000e+02,1.990000000000000000e+02,1.980000000000000000e+02,1.980000000000000000e+02,1.900000000000000000e+02,1.840000000000000000e+02,1.710000000000000000e+02,1.330000000000000000e+02,4.400000000000000000e+01,3.900000000000000000e+01,3.300000000000000000e+01,1.800000000000000000e+01,7.000000000000000000e+00,8.000000000000000000e+00,1.300000000000000000e+01,1.300000000000000000e+01,1.100000000000000000e+01,1.400000000000000000e+01,1.200000000000000000e+01,1.300000000000000000e+01,1.200000000000000000e+01,1.200000000000000000e+01,1.300000000000000000e+01,1.100000000000000000e+01,1.100000000000000000e+01,1.100000000000000000e+01,1.400000000000000000e+01,1.400000000000000000e+01),
(1.400000000000000000e+02,1.240000000000000000e+02,9.400000000000000000e+01,6.500000000000000000e+01,4.700000000000000000e+01,3.700000000000000000e+01,6.300000000000000000e+01,9.000000000000000000e+01,1.290000000000000000e+02,1.290000000000000000e+02,1.070000000000000000e+02,7.700000000000000000e+01,3.800000000000000000e+01,1.700000000000000000e+01,4.000000000000000000e+00,8.000000000000000000e+00,7.000000000000000000e+00,9.000000000000000000e+00,1.000000000000000000e+01,3.700000000000000000e+01,5.200000000000000000e+01,8.200000000000000000e+01,1.810000000000000000e+02,1.740000000000000000e+02,1.650000000000000000e+02,1.550000000000000000e+02,1.610000000000000000e+02,1.630000000000000000e+02,1.740000000000000000e+02,1.710000000000000000e+02,1.580000000000000000e+02,1.490000000000000000e+02,1.440000000000000000e+02,1.370000000000000000e+02,1.580000000000000000e+02,1.620000000000000000e+02,1.710000000000000000e+02,1.830000000000000000e+02,1.960000000000000000e+02,1.710000000000000000e+02,1.610000000000000000e+02,1.750000000000000000e+02,1.890000000000000000e+02,1.760000000000000000e+02,1.640000000000000000e+02,1.360000000000000000e+02,1.780000000000000000e+02,1.590000000000000000e+02,1.530000000000000000e+02,1.840000000000000000e+02,1.750000000000000000e+02,1.460000000000000000e+02,1.080000000000000000e+02,9.800000000000000000e+01,1.180000000000000000e+02,3.600000000000000000e+01,1.100000000000000000e+02,2.800000000000000000e+01,6.200000000000000000e+01,1.090000000000000000e+02,6.600000000000000000e+01,5.400000000000000000e+01,6.100000000000000000e+01,8.000000000000000000e+01,3.300000000000000000e+01,1.900000000000000000e+01,3.000000000000000000e+00,9.000000000000000000e+00,1.800000000000000000e+01,1.400000000000000000e+01,1.000000000000000000e+01,1.100000000000000000e+01,8.000000000000000000e+00,1.300000000000000000e+01,2.800000000000000000e+01,4.900000000000000000e+01,4.300000000000000000e+01,3.700000000000000000e+01,3.200000000000000000e+01,4.400000000000000000e+01,5.200000000000000000e+01,6.400000000000000000e+01,9.800000000000000000e+01,1.080000000000000000e+02,8.300000000000000000e+01,1.030000000000000000e+02,9.500000000000000000e+01,8.600000000000000000e+01,1.150000000000000000e+02,1.530000000000000000e+02,1.420000000000000000e+02,1.620000000000000000e+02,1.860000000000000000e+02,1.880000000000000000e+02,1.990000000000000000e+02,2.010000000000000000e+02,1.940000000000000000e+02,1.960000000000000000e+02,1.980000000000000000e+02,1.960000000000000000e+02,2.000000000000000000e+02,2.010000000000000000e+02,2.010000000000000000e+02,1.970000000000000000e+02,1.880000000000000000e+02,1.740000000000000000e+02,1.610000000000000000e+02,1.430000000000000000e+02,6.300000000000000000e+01,4.900000000000000000e+01,4.000000000000000000e+01,3.700000000000000000e+01,3.400000000000000000e+01,3.900000000000000000e+01,4.300000000000000000e+01,4.900000000000000000e+01,5.500000000000000000e+01,5.400000000000000000e+01,5.300000000000000000e+01,5.600000000000000000e+01,5.200000000000000000e+01,5.200000000000000000e+01,5.200000000000000000e+01,5.300000000000000000e+01,5.500000000000000000e+01,5.500000000000000000e+01,5.700000000000000000e+01,5.200000000000000000e+01),
(1.400000000000000000e+02,1.270000000000000000e+02,9.100000000000000000e+01,6.800000000000000000e+01,4.700000000000000000e+01,3.700000000000000000e+01,6.400000000000000000e+01,9.200000000000000000e+01,1.260000000000000000e+02,1.190000000000000000e+02,1.030000000000000000e+02,8.000000000000000000e+01,4.100000000000000000e+01,1.600000000000000000e+01,9.000000000000000000e+00,1.500000000000000000e+01,1.600000000000000000e+01,1.700000000000000000e+01,1.900000000000000000e+01,4.600000000000000000e+01,6.900000000000000000e+01,9.200000000000000000e+01,1.700000000000000000e+02,1.830000000000000000e+02,1.650000000000000000e+02,1.600000000000000000e+02,1.570000000000000000e+02,1.640000000000000000e+02,1.580000000000000000e+02,1.720000000000000000e+02,1.750000000000000000e+02,1.620000000000000000e+02,1.610000000000000000e+02,1.700000000000000000e+02,1.560000000000000000e+02,1.550000000000000000e+02,1.510000000000000000e+02,1.800000000000000000e+02,1.900000000000000000e+02,1.860000000000000000e+02,1.610000000000000000e+02,1.890000000000000000e+02,1.890000000000000000e+02,1.790000000000000000e+02,1.730000000000000000e+02,1.680000000000000000e+02,1.730000000000000000e+02,1.630000000000000000e+02,1.600000000000000000e+02,1.640000000000000000e+02,1.700000000000000000e+02,1.510000000000000000e+02,1.380000000000000000e+02,1.040000000000000000e+02,4.300000000000000000e+01,4.200000000000000000e+01,4.200000000000000000e+01,4.200000000000000000e+01,2.100000000000000000e+01,9.900000000000000000e+01,4.500000000000000000e+01,7.400000000000000000e+01,1.170000000000000000e+02,6.800000000000000000e+01,3.400000000000000000e+01,1.200000000000000000e+01,8.000000000000000000e+00,7.000000000000000000e+00,9.000000000000000000e+00,1.400000000000000000e+01,8.000000000000000000e+00,1.200000000000000000e+01,1.200000000000000000e+01,1.800000000000000000e+01,2.400000000000000000e+01,3.000000000000000000e+01,4.000000000000000000e+01,2.000000000000000000e+01,3.300000000000000000e+01,3.900000000000000000e+01,3.700000000000000000e+01,5.000000000000000000e+01,5.600000000000000000e+01,7.800000000000000000e+01,8.100000000000000000e+01,6.800000000000000000e+01,8.000000000000000000e+01,1.050000000000000000e+02,1.290000000000000000e+02,1.560000000000000000e+02,1.590000000000000000e+02,1.150000000000000000e+02,1.490000000000000000e+02,1.530000000000000000e+02,1.510000000000000000e+02,1.640000000000000000e+02,1.860000000000000000e+02,1.890000000000000000e+02,1.950000000000000000e+02,1.960000000000000000e+02,1.990000000000000000e+02,2.050000000000000000e+02,1.980000000000000000e+02,1.850000000000000000e+02,1.800000000000000000e+02,1.700000000000000000e+02,1.510000000000000000e+02,1.340000000000000000e+02,9.800000000000000000e+01,9.800000000000000000e+01,8.200000000000000000e+01,8.000000000000000000e+01,8.100000000000000000e+01,8.300000000000000000e+01,8.200000000000000000e+01,9.400000000000000000e+01,1.050000000000000000e+02,1.060000000000000000e+02,1.090000000000000000e+02,1.100000000000000000e+02,1.030000000000000000e+02,1.060000000000000000e+02,1.030000000000000000e+02,1.040000000000000000e+02,1.060000000000000000e+02,1.060000000000000000e+02,1.060000000000000000e+02,1.020000000000000000e+02),
(1.440000000000000000e+02,1.280000000000000000e+02,9.700000000000000000e+01,7.000000000000000000e+01,5.200000000000000000e+01,3.700000000000000000e+01,6.100000000000000000e+01,9.100000000000000000e+01,1.230000000000000000e+02,1.200000000000000000e+02,1.040000000000000000e+02,8.200000000000000000e+01,5.400000000000000000e+01,3.100000000000000000e+01,2.600000000000000000e+01,3.100000000000000000e+01,3.600000000000000000e+01,4.000000000000000000e+01,4.200000000000000000e+01,8.000000000000000000e+01,8.000000000000000000e+01,1.210000000000000000e+02,1.310000000000000000e+02,1.670000000000000000e+02,1.610000000000000000e+02,1.830000000000000000e+02,1.900000000000000000e+02,1.810000000000000000e+02,1.690000000000000000e+02,1.830000000000000000e+02,1.900000000000000000e+02,1.890000000000000000e+02,1.940000000000000000e+02,1.960000000000000000e+02,1.980000000000000000e+02,2.010000000000000000e+02,1.980000000000000000e+02,1.920000000000000000e+02,1.950000000000000000e+02,1.870000000000000000e+02,1.710000000000000000e+02,1.900000000000000000e+02,1.940000000000000000e+02,1.690000000000000000e+02,1.670000000000000000e+02,2.010000000000000000e+02,1.760000000000000000e+02,1.960000000000000000e+02,1.570000000000000000e+02,1.790000000000000000e+02,1.540000000000000000e+02,1.480000000000000000e+02,9.200000000000000000e+01,7.600000000000000000e+01,3.500000000000000000e+01,5.900000000000000000e+01,6.200000000000000000e+01,3.400000000000000000e+01,4.400000000000000000e+01,3.700000000000000000e+01,9.500000000000000000e+01,1.230000000000000000e+02,7.000000000000000000e+01,1.210000000000000000e+02,5.200000000000000000e+01,5.000000000000000000e+00,2.900000000000000000e+01,3.000000000000000000e+01,4.100000000000000000e+01,1.400000000000000000e+01,6.000000000000000000e+00,6.000000000000000000e+00,1.600000000000000000e+01,1.200000000000000000e+01,2.200000000000000000e+01,1.400000000000000000e+01,2.200000000000000000e+01,1.900000000000000000e+01,1.600000000000000000e+01,2.500000000000000000e+01,5.000000000000000000e+01,2.300000000000000000e+01,1.500000000000000000e+01,5.400000000000000000e+01,4.400000000000000000e+01,3.900000000000000000e+01,8.900000000000000000e+01,1.340000000000000000e+02,1.540000000000000000e+02,1.770000000000000000e+02,1.740000000000000000e+02,1.350000000000000000e+02,1.640000000000000000e+02,1.650000000000000000e+02,1.730000000000000000e+02,1.830000000000000000e+02,1.800000000000000000e+02,1.830000000000000000e+02,1.940000000000000000e+02,1.970000000000000000e+02,1.990000000000000000e+02,1.970000000000000000e+02,1.940000000000000000e+02,1.770000000000000000e+02,1.710000000000000000e+02,1.550000000000000000e+02,1.640000000000000000e+02,1.520000000000000000e+02,1.440000000000000000e+02,1.430000000000000000e+02,1.250000000000000000e+02,1.200000000000000000e+02,1.190000000000000000e+02,1.220000000000000000e+02,1.190000000000000000e+02,1.340000000000000000e+02,1.440000000000000000e+02,1.510000000000000000e+02,1.480000000000000000e+02,1.480000000000000000e+02,1.440000000000000000e+02,1.460000000000000000e+02,1.480000000000000000e+02,1.420000000000000000e+02,1.470000000000000000e+02,1.480000000000000000e+02,1.480000000000000000e+02,1.470000000000000000e+02),
(1.410000000000000000e+02,1.280000000000000000e+02,9.700000000000000000e+01,6.900000000000000000e+01,4.900000000000000000e+01,3.700000000000000000e+01,6.900000000000000000e+01,9.300000000000000000e+01,1.270000000000000000e+02,1.250000000000000000e+02,1.170000000000000000e+02,9.300000000000000000e+01,7.200000000000000000e+01,5.100000000000000000e+01,5.900000000000000000e+01,6.600000000000000000e+01,7.500000000000000000e+01,7.400000000000000000e+01,7.000000000000000000e+01,8.100000000000000000e+01,9.600000000000000000e+01,1.460000000000000000e+02,1.040000000000000000e+02,1.380000000000000000e+02,1.870000000000000000e+02,2.050000000000000000e+02,1.900000000000000000e+02,1.920000000000000000e+02,1.790000000000000000e+02,1.940000000000000000e+02,1.950000000000000000e+02,1.950000000000000000e+02,1.940000000000000000e+02,1.930000000000000000e+02,1.870000000000000000e+02,1.910000000000000000e+02,1.950000000000000000e+02,1.750000000000000000e+02,1.650000000000000000e+02,1.550000000000000000e+02,1.860000000000000000e+02,1.960000000000000000e+02,1.960000000000000000e+02,1.880000000000000000e+02,1.820000000000000000e+02,2.000000000000000000e+02,1.940000000000000000e+02,2.010000000000000000e+02,1.990000000000000000e+02,1.850000000000000000e+02,1.560000000000000000e+02,1.330000000000000000e+02,1.070000000000000000e+02,9.000000000000000000e+01,4.300000000000000000e+01,4.800000000000000000e+01,1.500000000000000000e+01,5.000000000000000000e+01,2.300000000000000000e+01,2.700000000000000000e+01,5.400000000000000000e+01,8.800000000000000000e+01,5.600000000000000000e+01,8.000000000000000000e+01,6.300000000000000000e+01,1.100000000000000000e+01,1.600000000000000000e+01,9.900000000000000000e+01,7.100000000000000000e+01,4.900000000000000000e+01,1.800000000000000000e+01,9.000000000000000000e+00,4.700000000000000000e+01,9.000000000000000000e+00,2.000000000000000000e+01,5.100000000000000000e+01,1.100000000000000000e+01,5.400000000000000000e+01,2.000000000000000000e+01,6.000000000000000000e+00,2.100000000000000000e+01,3.500000000000000000e+01,2.500000000000000000e+01,2.000000000000000000e+01,4.000000000000000000e+01,3.300000000000000000e+01,8.300000000000000000e+01,1.140000000000000000e+02,1.460000000000000000e+02,2.000000000000000000e+02,1.530000000000000000e+02,1.580000000000000000e+02,1.850000000000000000e+02,1.740000000000000000e+02,1.800000000000000000e+02,1.670000000000000000e+02,1.730000000000000000e+02,1.880000000000000000e+02,1.940000000000000000e+02,1.990000000000000000e+02,1.980000000000000000e+02,1.860000000000000000e+02,1.790000000000000000e+02,1.740000000000000000e+02,1.750000000000000000e+02,1.590000000000000000e+02,1.730000000000000000e+02,1.790000000000000000e+02,1.820000000000000000e+02,1.770000000000000000e+02,1.600000000000000000e+02,1.560000000000000000e+02,1.530000000000000000e+02,1.560000000000000000e+02,1.540000000000000000e+02,1.630000000000000000e+02,1.770000000000000000e+02,1.770000000000000000e+02,1.730000000000000000e+02,1.760000000000000000e+02,1.720000000000000000e+02,1.710000000000000000e+02,1.750000000000000000e+02,1.770000000000000000e+02,1.770000000000000000e+02,1.730000000000000000e+02,1.760000000000000000e+02,1.780000000000000000e+02),
(1.470000000000000000e+02,1.320000000000000000e+02,1.000000000000000000e+02,6.700000000000000000e+01,4.700000000000000000e+01,3.900000000000000000e+01,6.500000000000000000e+01,9.600000000000000000e+01,1.350000000000000000e+02,1.290000000000000000e+02,1.110000000000000000e+02,9.700000000000000000e+01,8.500000000000000000e+01,7.300000000000000000e+01,7.600000000000000000e+01,9.800000000000000000e+01,1.040000000000000000e+02,1.040000000000000000e+02,1.000000000000000000e+02,8.200000000000000000e+01,1.030000000000000000e+02,1.590000000000000000e+02,1.300000000000000000e+02,1.050000000000000000e+02,2.030000000000000000e+02,1.880000000000000000e+02,1.510000000000000000e+02,1.820000000000000000e+02,1.690000000000000000e+02,1.610000000000000000e+02,1.670000000000000000e+02,1.840000000000000000e+02,1.860000000000000000e+02,1.860000000000000000e+02,1.870000000000000000e+02,1.980000000000000000e+02,1.880000000000000000e+02,1.890000000000000000e+02,1.590000000000000000e+02,1.620000000000000000e+02,1.840000000000000000e+02,1.970000000000000000e+02,2.020000000000000000e+02,1.900000000000000000e+02,1.750000000000000000e+02,1.940000000000000000e+02,2.010000000000000000e+02,1.870000000000000000e+02,1.910000000000000000e+02,1.780000000000000000e+02,1.200000000000000000e+02,6.300000000000000000e+01,4.500000000000000000e+01,1.300000000000000000e+01,3.000000000000000000e+01,9.800000000000000000e+01,8.000000000000000000e+01,6.300000000000000000e+01,2.400000000000000000e+01,3.000000000000000000e+01,8.000000000000000000e+00,3.000000000000000000e+01,2.500000000000000000e+01,8.600000000000000000e+01,7.700000000000000000e+01,1.700000000000000000e+01,1.000000000000000000e+01,8.000000000000000000e+01,1.210000000000000000e+02,5.800000000000000000e+01,2.000000000000000000e+01,4.000000000000000000e+00,5.400000000000000000e+01,6.000000000000000000e+00,6.000000000000000000e+00,2.800000000000000000e+01,3.600000000000000000e+01,2.400000000000000000e+01,8.000000000000000000e+01,6.000000000000000000e+00,9.000000000000000000e+00,2.800000000000000000e+01,2.100000000000000000e+01,3.000000000000000000e+01,3.000000000000000000e+01,5.800000000000000000e+01,1.080000000000000000e+02,8.200000000000000000e+01,1.510000000000000000e+02,1.960000000000000000e+02,1.660000000000000000e+02,2.000000000000000000e+02,1.980000000000000000e+02,1.900000000000000000e+02,1.800000000000000000e+02,1.740000000000000000e+02,1.750000000000000000e+02,1.800000000000000000e+02,1.920000000000000000e+02,1.990000000000000000e+02,1.850000000000000000e+02,1.760000000000000000e+02,1.770000000000000000e+02,1.930000000000000000e+02,1.800000000000000000e+02,1.680000000000000000e+02,1.780000000000000000e+02,1.870000000000000000e+02,1.890000000000000000e+02,1.870000000000000000e+02,1.740000000000000000e+02,1.700000000000000000e+02,1.660000000000000000e+02,1.680000000000000000e+02,1.690000000000000000e+02,1.790000000000000000e+02,1.880000000000000000e+02,1.850000000000000000e+02,1.870000000000000000e+02,1.860000000000000000e+02,1.860000000000000000e+02,1.860000000000000000e+02,1.840000000000000000e+02,1.840000000000000000e+02,1.820000000000000000e+02,1.850000000000000000e+02,1.830000000000000000e+02,1.820000000000000000e+02),
(1.430000000000000000e+02,1.270000000000000000e+02,9.300000000000000000e+01,6.800000000000000000e+01,4.400000000000000000e+01,3.600000000000000000e+01,6.700000000000000000e+01,1.000000000000000000e+02,1.320000000000000000e+02,1.230000000000000000e+02,1.200000000000000000e+02,1.110000000000000000e+02,9.800000000000000000e+01,9.600000000000000000e+01,1.020000000000000000e+02,1.190000000000000000e+02,1.290000000000000000e+02,1.230000000000000000e+02,9.500000000000000000e+01,8.000000000000000000e+01,9.900000000000000000e+01,1.790000000000000000e+02,1.750000000000000000e+02,1.120000000000000000e+02,1.980000000000000000e+02,1.690000000000000000e+02,1.270000000000000000e+02,1.760000000000000000e+02,1.440000000000000000e+02,1.540000000000000000e+02,1.510000000000000000e+02,1.710000000000000000e+02,1.820000000000000000e+02,1.900000000000000000e+02,1.890000000000000000e+02,2.020000000000000000e+02,1.830000000000000000e+02,1.880000000000000000e+02,1.870000000000000000e+02,1.730000000000000000e+02,1.920000000000000000e+02,2.020000000000000000e+02,1.900000000000000000e+02,1.940000000000000000e+02,1.920000000000000000e+02,1.950000000000000000e+02,1.820000000000000000e+02,1.550000000000000000e+02,1.590000000000000000e+02,1.550000000000000000e+02,1.620000000000000000e+02,2.400000000000000000e+01,4.300000000000000000e+01,2.800000000000000000e+01,7.100000000000000000e+01,9.500000000000000000e+01,1.590000000000000000e+02,8.500000000000000000e+01,1.380000000000000000e+02,3.700000000000000000e+01,1.000000000000000000e+01,1.430000000000000000e+02,1.040000000000000000e+02,5.400000000000000000e+01,7.500000000000000000e+01,1.700000000000000000e+01,2.600000000000000000e+01,5.000000000000000000e+01,6.900000000000000000e+01,5.400000000000000000e+01,1.300000000000000000e+02,2.200000000000000000e+01,1.500000000000000000e+01,1.000000000000000000e+01,2.900000000000000000e+01,1.500000000000000000e+01,3.300000000000000000e+01,6.000000000000000000e+00,5.600000000000000000e+01,5.100000000000000000e+01,4.000000000000000000e+00,1.200000000000000000e+01,4.500000000000000000e+01,1.200000000000000000e+01,1.700000000000000000e+01,6.300000000000000000e+01,7.600000000000000000e+01,8.600000000000000000e+01,1.200000000000000000e+02,1.530000000000000000e+02,1.850000000000000000e+02,1.970000000000000000e+02,2.060000000000000000e+02,2.000000000000000000e+02,1.900000000000000000e+02,1.810000000000000000e+02,1.800000000000000000e+02,1.870000000000000000e+02,1.920000000000000000e+02,1.700000000000000000e+02,1.700000000000000000e+02,1.860000000000000000e+02,1.910000000000000000e+02,1.930000000000000000e+02,1.790000000000000000e+02,1.740000000000000000e+02,1.810000000000000000e+02,1.840000000000000000e+02,1.880000000000000000e+02,1.860000000000000000e+02,1.760000000000000000e+02,1.630000000000000000e+02,1.630000000000000000e+02,1.680000000000000000e+02,1.660000000000000000e+02,1.760000000000000000e+02,1.850000000000000000e+02,1.790000000000000000e+02,1.810000000000000000e+02,1.830000000000000000e+02,1.830000000000000000e+02,1.860000000000000000e+02,1.860000000000000000e+02,1.860000000000000000e+02,1.850000000000000000e+02,1.850000000000000000e+02,1.860000000000000000e+02,1.850000000000000000e+02),
(1.460000000000000000e+02,1.250000000000000000e+02,9.700000000000000000e+01,6.500000000000000000e+01,4.400000000000000000e+01,4.100000000000000000e+01,7.300000000000000000e+01,9.900000000000000000e+01,1.300000000000000000e+02,1.300000000000000000e+02,1.220000000000000000e+02,1.120000000000000000e+02,1.040000000000000000e+02,1.050000000000000000e+02,1.140000000000000000e+02,1.230000000000000000e+02,1.270000000000000000e+02,1.300000000000000000e+02,1.030000000000000000e+02,7.300000000000000000e+01,1.090000000000000000e+02,1.750000000000000000e+02,2.040000000000000000e+02,1.980000000000000000e+02,1.750000000000000000e+02,1.440000000000000000e+02,1.290000000000000000e+02,1.620000000000000000e+02,1.260000000000000000e+02,1.270000000000000000e+02,1.710000000000000000e+02,1.890000000000000000e+02,1.990000000000000000e+02,2.090000000000000000e+02,2.060000000000000000e+02,2.090000000000000000e+02,1.980000000000000000e+02,1.890000000000000000e+02,1.910000000000000000e+02,1.950000000000000000e+02,1.990000000000000000e+02,1.890000000000000000e+02,1.940000000000000000e+02,1.660000000000000000e+02,1.880000000000000000e+02,1.680000000000000000e+02,1.260000000000000000e+02,1.270000000000000000e+02,8.800000000000000000e+01,1.060000000000000000e+02,1.400000000000000000e+02,4.300000000000000000e+01,1.010000000000000000e+02,5.800000000000000000e+01,1.200000000000000000e+02,1.530000000000000000e+02,5.300000000000000000e+01,1.530000000000000000e+02,1.420000000000000000e+02,6.500000000000000000e+01,7.300000000000000000e+01,1.440000000000000000e+02,1.260000000000000000e+02,1.230000000000000000e+02,9.700000000000000000e+01,3.800000000000000000e+01,3.600000000000000000e+01,2.600000000000000000e+01,1.700000000000000000e+01,3.700000000000000000e+01,1.310000000000000000e+02,9.700000000000000000e+01,2.700000000000000000e+01,3.800000000000000000e+01,2.100000000000000000e+01,1.100000000000000000e+01,1.800000000000000000e+01,1.300000000000000000e+01,1.360000000000000000e+02,3.200000000000000000e+01,1.100000000000000000e+01,1.000000000000000000e+00,7.000000000000000000e+00,3.600000000000000000e+01,5.500000000000000000e+01,3.900000000000000000e+01,4.100000000000000000e+01,5.900000000000000000e+01,8.300000000000000000e+01,8.200000000000000000e+01,1.810000000000000000e+02,1.960000000000000000e+02,2.060000000000000000e+02,1.970000000000000000e+02,2.070000000000000000e+02,2.070000000000000000e+02,2.070000000000000000e+02,2.020000000000000000e+02,1.980000000000000000e+02,1.940000000000000000e+02,2.020000000000000000e+02,2.040000000000000000e+02,2.000000000000000000e+02,1.990000000000000000e+02,1.920000000000000000e+02,1.890000000000000000e+02,1.770000000000000000e+02,1.790000000000000000e+02,1.810000000000000000e+02,1.800000000000000000e+02,1.680000000000000000e+02,1.620000000000000000e+02,1.560000000000000000e+02,1.600000000000000000e+02,1.530000000000000000e+02,1.660000000000000000e+02,1.720000000000000000e+02,1.690000000000000000e+02,1.760000000000000000e+02,1.810000000000000000e+02,1.800000000000000000e+02,1.850000000000000000e+02,1.860000000000000000e+02,1.860000000000000000e+02,1.870000000000000000e+02,1.870000000000000000e+02,1.860000000000000000e+02,1.870000000000000000e+02),
(1.430000000000000000e+02,1.260000000000000000e+02,9.800000000000000000e+01,6.100000000000000000e+01,4.400000000000000000e+01,4.000000000000000000e+01,7.500000000000000000e+01,9.900000000000000000e+01,1.310000000000000000e+02,1.290000000000000000e+02,1.220000000000000000e+02,1.120000000000000000e+02,1.090000000000000000e+02,1.030000000000000000e+02,1.060000000000000000e+02,1.120000000000000000e+02,1.160000000000000000e+02,1.090000000000000000e+02,9.500000000000000000e+01,7.200000000000000000e+01,9.400000000000000000e+01,1.840000000000000000e+02,2.090000000000000000e+02,2.030000000000000000e+02,1.680000000000000000e+02,1.340000000000000000e+02,1.280000000000000000e+02,1.480000000000000000e+02,1.030000000000000000e+02,1.440000000000000000e+02,1.890000000000000000e+02,1.980000000000000000e+02,2.100000000000000000e+02,2.110000000000000000e+02,2.110000000000000000e+02,2.110000000000000000e+02,2.060000000000000000e+02,2.070000000000000000e+02,2.070000000000000000e+02,2.000000000000000000e+02,1.890000000000000000e+02,1.870000000000000000e+02,1.460000000000000000e+02,1.810000000000000000e+02,1.380000000000000000e+02,1.460000000000000000e+02,1.160000000000000000e+02,1.430000000000000000e+02,6.400000000000000000e+01,8.100000000000000000e+01,1.570000000000000000e+02,5.400000000000000000e+01,1.620000000000000000e+02,1.400000000000000000e+02,1.000000000000000000e+02,1.550000000000000000e+02,9.900000000000000000e+01,6.300000000000000000e+01,4.900000000000000000e+01,9.100000000000000000e+01,9.600000000000000000e+01,1.260000000000000000e+02,9.800000000000000000e+01,1.440000000000000000e+02,6.200000000000000000e+01,6.600000000000000000e+01,2.100000000000000000e+01,7.000000000000000000e+00,1.000000000000000000e+01,5.800000000000000000e+01,1.850000000000000000e+02,1.010000000000000000e+02,7.300000000000000000e+01,5.700000000000000000e+01,1.700000000000000000e+01,1.600000000000000000e+01,2.500000000000000000e+01,3.900000000000000000e+01,2.010000000000000000e+02,9.800000000000000000e+01,1.300000000000000000e+01,1.000000000000000000e+00,9.000000000000000000e+00,7.400000000000000000e+01,8.500000000000000000e+01,6.200000000000000000e+01,2.100000000000000000e+01,5.900000000000000000e+01,5.700000000000000000e+01,8.500000000000000000e+01,1.330000000000000000e+02,1.970000000000000000e+02,1.790000000000000000e+02,2.000000000000000000e+02,2.060000000000000000e+02,2.050000000000000000e+02,2.030000000000000000e+02,2.000000000000000000e+02,2.070000000000000000e+02,2.020000000000000000e+02,2.050000000000000000e+02,2.060000000000000000e+02,2.070000000000000000e+02,2.030000000000000000e+02,2.000000000000000000e+02,1.840000000000000000e+02,1.770000000000000000e+02,1.760000000000000000e+02,1.780000000000000000e+02,1.770000000000000000e+02,1.620000000000000000e+02,1.620000000000000000e+02,1.610000000000000000e+02,1.580000000000000000e+02,1.630000000000000000e+02,1.710000000000000000e+02,1.750000000000000000e+02,1.720000000000000000e+02,1.680000000000000000e+02,1.680000000000000000e+02,1.700000000000000000e+02,1.770000000000000000e+02,1.820000000000000000e+02,1.790000000000000000e+02,1.800000000000000000e+02,1.820000000000000000e+02,1.840000000000000000e+02,1.800000000000000000e+02),
(1.400000000000000000e+02,1.220000000000000000e+02,8.400000000000000000e+01,6.200000000000000000e+01,4.100000000000000000e+01,4.000000000000000000e+01,7.400000000000000000e+01,1.040000000000000000e+02,1.440000000000000000e+02,1.310000000000000000e+02,1.240000000000000000e+02,1.130000000000000000e+02,1.030000000000000000e+02,1.000000000000000000e+02,1.020000000000000000e+02,1.070000000000000000e+02,9.700000000000000000e+01,1.000000000000000000e+02,7.300000000000000000e+01,6.400000000000000000e+01,9.300000000000000000e+01,1.830000000000000000e+02,2.060000000000000000e+02,2.040000000000000000e+02,1.540000000000000000e+02,1.390000000000000000e+02,1.210000000000000000e+02,1.550000000000000000e+02,8.800000000000000000e+01,1.130000000000000000e+02,1.690000000000000000e+02,1.820000000000000000e+02,1.980000000000000000e+02,1.990000000000000000e+02,2.070000000000000000e+02,2.080000000000000000e+02,2.080000000000000000e+02,2.010000000000000000e+02,2.070000000000000000e+02,2.040000000000000000e+02,1.680000000000000000e+02,1.830000000000000000e+02,1.380000000000000000e+02,1.710000000000000000e+02,1.310000000000000000e+02,1.190000000000000000e+02,1.420000000000000000e+02,8.600000000000000000e+01,8.300000000000000000e+01,8.900000000000000000e+01,1.380000000000000000e+02,1.050000000000000000e+02,1.160000000000000000e+02,1.370000000000000000e+02,1.160000000000000000e+02,1.340000000000000000e+02,1.390000000000000000e+02,1.300000000000000000e+02,4.900000000000000000e+01,1.280000000000000000e+02,1.150000000000000000e+02,1.150000000000000000e+02,9.900000000000000000e+01,1.120000000000000000e+02,1.050000000000000000e+02,2.100000000000000000e+01,1.000000000000000000e+00,1.100000000000000000e+01,1.200000000000000000e+01,2.200000000000000000e+01,3.300000000000000000e+01,9.700000000000000000e+01,1.030000000000000000e+02,4.400000000000000000e+01,3.300000000000000000e+01,2.300000000000000000e+01,8.800000000000000000e+01,4.100000000000000000e+01,1.860000000000000000e+02,7.100000000000000000e+01,3.500000000000000000e+01,1.000000000000000000e+00,7.000000000000000000e+00,4.700000000000000000e+01,4.600000000000000000e+01,3.300000000000000000e+01,4.400000000000000000e+01,6.900000000000000000e+01,5.000000000000000000e+01,4.800000000000000000e+01,1.160000000000000000e+02,1.740000000000000000e+02,1.790000000000000000e+02,2.000000000000000000e+02,2.040000000000000000e+02,2.050000000000000000e+02,2.030000000000000000e+02,2.040000000000000000e+02,2.060000000000000000e+02,2.030000000000000000e+02,2.050000000000000000e+02,2.080000000000000000e+02,2.080000000000000000e+02,2.000000000000000000e+02,1.840000000000000000e+02,1.490000000000000000e+02,1.630000000000000000e+02,1.660000000000000000e+02,1.680000000000000000e+02,1.680000000000000000e+02,1.670000000000000000e+02,1.580000000000000000e+02,1.530000000000000000e+02,1.530000000000000000e+02,1.630000000000000000e+02,1.690000000000000000e+02,1.680000000000000000e+02,1.670000000000000000e+02,1.690000000000000000e+02,1.680000000000000000e+02,1.740000000000000000e+02,1.770000000000000000e+02,1.840000000000000000e+02,1.780000000000000000e+02,1.660000000000000000e+02,1.670000000000000000e+02,1.640000000000000000e+02,1.630000000000000000e+02),
(1.410000000000000000e+02,1.180000000000000000e+02,8.700000000000000000e+01,5.900000000000000000e+01,4.100000000000000000e+01,3.600000000000000000e+01,6.900000000000000000e+01,1.030000000000000000e+02,1.400000000000000000e+02,1.320000000000000000e+02,1.260000000000000000e+02,1.130000000000000000e+02,1.040000000000000000e+02,9.300000000000000000e+01,9.600000000000000000e+01,9.700000000000000000e+01,8.600000000000000000e+01,7.500000000000000000e+01,7.000000000000000000e+01,5.000000000000000000e+01,8.800000000000000000e+01,1.750000000000000000e+02,2.010000000000000000e+02,1.970000000000000000e+02,1.380000000000000000e+02,1.190000000000000000e+02,1.340000000000000000e+02,1.680000000000000000e+02,1.170000000000000000e+02,1.340000000000000000e+02,1.640000000000000000e+02,1.730000000000000000e+02,1.830000000000000000e+02,1.590000000000000000e+02,2.010000000000000000e+02,2.050000000000000000e+02,1.980000000000000000e+02,2.020000000000000000e+02,2.090000000000000000e+02,1.900000000000000000e+02,1.370000000000000000e+02,1.740000000000000000e+02,1.440000000000000000e+02,1.430000000000000000e+02,1.780000000000000000e+02,1.390000000000000000e+02,1.480000000000000000e+02,9.600000000000000000e+01,9.400000000000000000e+01,1.020000000000000000e+02,1.340000000000000000e+02,1.420000000000000000e+02,1.070000000000000000e+02,1.200000000000000000e+02,1.500000000000000000e+02,1.220000000000000000e+02,1.170000000000000000e+02,6.000000000000000000e+01,5.000000000000000000e+01,2.300000000000000000e+01,6.600000000000000000e+01,3.400000000000000000e+01,1.250000000000000000e+02,1.570000000000000000e+02,9.100000000000000000e+01,3.900000000000000000e+01,5.000000000000000000e+00,2.200000000000000000e+01,2.000000000000000000e+01,6.100000000000000000e+01,6.300000000000000000e+01,8.900000000000000000e+01,1.210000000000000000e+02,1.700000000000000000e+02,4.300000000000000000e+01,1.800000000000000000e+01,6.500000000000000000e+01,4.500000000000000000e+01,1.680000000000000000e+02,8.900000000000000000e+01,2.600000000000000000e+01,8.000000000000000000e+00,1.200000000000000000e+01,9.000000000000000000e+00,7.300000000000000000e+01,6.300000000000000000e+01,9.700000000000000000e+01,8.000000000000000000e+01,6.900000000000000000e+01,4.900000000000000000e+01,1.520000000000000000e+02,1.110000000000000000e+02,1.800000000000000000e+02,1.990000000000000000e+02,1.920000000000000000e+02,2.030000000000000000e+02,2.060000000000000000e+02,2.040000000000000000e+02,2.060000000000000000e+02,2.030000000000000000e+02,2.080000000000000000e+02,2.080000000000000000e+02,2.030000000000000000e+02,1.670000000000000000e+02,8.500000000000000000e+01,1.220000000000000000e+02,1.490000000000000000e+02,1.600000000000000000e+02,1.650000000000000000e+02,1.740000000000000000e+02,1.640000000000000000e+02,1.590000000000000000e+02,1.470000000000000000e+02,1.470000000000000000e+02,1.560000000000000000e+02,1.680000000000000000e+02,1.650000000000000000e+02,1.610000000000000000e+02,1.600000000000000000e+02,1.590000000000000000e+02,1.670000000000000000e+02,1.700000000000000000e+02,1.660000000000000000e+02,1.570000000000000000e+02,1.460000000000000000e+02,1.380000000000000000e+02,1.340000000000000000e+02,1.280000000000000000e+02),
(1.350000000000000000e+02,1.180000000000000000e+02,8.400000000000000000e+01,6.100000000000000000e+01,4.000000000000000000e+01,3.800000000000000000e+01,7.700000000000000000e+01,1.020000000000000000e+02,1.340000000000000000e+02,1.290000000000000000e+02,1.310000000000000000e+02,1.140000000000000000e+02,1.080000000000000000e+02,9.400000000000000000e+01,9.400000000000000000e+01,9.600000000000000000e+01,8.600000000000000000e+01,8.100000000000000000e+01,8.000000000000000000e+01,5.500000000000000000e+01,7.900000000000000000e+01,1.070000000000000000e+02,1.690000000000000000e+02,1.840000000000000000e+02,1.230000000000000000e+02,8.200000000000000000e+01,1.410000000000000000e+02,1.770000000000000000e+02,1.340000000000000000e+02,1.420000000000000000e+02,1.320000000000000000e+02,1.470000000000000000e+02,1.670000000000000000e+02,1.900000000000000000e+02,1.970000000000000000e+02,2.040000000000000000e+02,1.720000000000000000e+02,1.880000000000000000e+02,1.820000000000000000e+02,1.560000000000000000e+02,1.390000000000000000e+02,1.550000000000000000e+02,1.530000000000000000e+02,1.380000000000000000e+02,1.910000000000000000e+02,1.030000000000000000e+02,1.200000000000000000e+02,1.280000000000000000e+02,1.030000000000000000e+02,1.030000000000000000e+02,1.050000000000000000e+02,1.540000000000000000e+02,1.450000000000000000e+02,1.720000000000000000e+02,1.010000000000000000e+02,1.150000000000000000e+02,5.600000000000000000e+01,4.100000000000000000e+01,2.700000000000000000e+01,1.000000000000000000e+01,2.600000000000000000e+01,1.000000000000000000e+02,9.200000000000000000e+01,1.320000000000000000e+02,7.800000000000000000e+01,2.300000000000000000e+01,8.400000000000000000e+01,1.310000000000000000e+02,1.060000000000000000e+02,8.400000000000000000e+01,3.600000000000000000e+01,7.600000000000000000e+01,1.180000000000000000e+02,1.760000000000000000e+02,2.800000000000000000e+01,2.300000000000000000e+01,3.200000000000000000e+01,1.800000000000000000e+01,1.590000000000000000e+02,1.000000000000000000e+02,1.700000000000000000e+01,2.600000000000000000e+01,6.000000000000000000e+00,3.600000000000000000e+01,8.500000000000000000e+01,6.800000000000000000e+01,6.600000000000000000e+01,6.100000000000000000e+01,9.900000000000000000e+01,1.590000000000000000e+02,8.500000000000000000e+01,1.360000000000000000e+02,1.670000000000000000e+02,1.850000000000000000e+02,1.860000000000000000e+02,2.010000000000000000e+02,2.080000000000000000e+02,2.040000000000000000e+02,2.030000000000000000e+02,1.850000000000000000e+02,1.900000000000000000e+02,1.960000000000000000e+02,1.940000000000000000e+02,1.600000000000000000e+02,9.200000000000000000e+01,1.270000000000000000e+02,1.430000000000000000e+02,1.540000000000000000e+02,1.650000000000000000e+02,1.700000000000000000e+02,1.670000000000000000e+02,1.580000000000000000e+02,1.530000000000000000e+02,1.520000000000000000e+02,1.530000000000000000e+02,1.590000000000000000e+02,1.640000000000000000e+02,1.530000000000000000e+02,1.530000000000000000e+02,1.600000000000000000e+02,1.530000000000000000e+02,1.490000000000000000e+02,1.420000000000000000e+02,1.290000000000000000e+02,1.070000000000000000e+02,1.010000000000000000e+02,8.500000000000000000e+01,8.500000000000000000e+01),
(1.380000000000000000e+02,1.240000000000000000e+02,9.000000000000000000e+01,6.100000000000000000e+01,3.800000000000000000e+01,3.700000000000000000e+01,7.100000000000000000e+01,1.020000000000000000e+02,1.340000000000000000e+02,1.270000000000000000e+02,1.250000000000000000e+02,1.130000000000000000e+02,1.040000000000000000e+02,9.500000000000000000e+01,9.400000000000000000e+01,9.200000000000000000e+01,8.200000000000000000e+01,7.600000000000000000e+01,7.800000000000000000e+01,5.100000000000000000e+01,5.700000000000000000e+01,1.120000000000000000e+02,9.400000000000000000e+01,1.620000000000000000e+02,1.290000000000000000e+02,8.700000000000000000e+01,8.900000000000000000e+01,1.770000000000000000e+02,1.710000000000000000e+02,1.590000000000000000e+02,1.760000000000000000e+02,1.920000000000000000e+02,1.990000000000000000e+02,2.020000000000000000e+02,1.940000000000000000e+02,2.060000000000000000e+02,2.010000000000000000e+02,1.960000000000000000e+02,1.060000000000000000e+02,1.780000000000000000e+02,1.550000000000000000e+02,1.140000000000000000e+02,1.480000000000000000e+02,1.420000000000000000e+02,1.740000000000000000e+02,1.420000000000000000e+02,1.370000000000000000e+02,1.340000000000000000e+02,1.190000000000000000e+02,1.080000000000000000e+02,1.550000000000000000e+02,9.800000000000000000e+01,1.000000000000000000e+02,1.280000000000000000e+02,1.620000000000000000e+02,4.500000000000000000e+01,5.900000000000000000e+01,7.400000000000000000e+01,1.300000000000000000e+02,7.500000000000000000e+01,3.900000000000000000e+01,7.200000000000000000e+01,5.200000000000000000e+01,8.800000000000000000e+01,2.400000000000000000e+01,2.000000000000000000e+01,1.220000000000000000e+02,1.270000000000000000e+02,1.480000000000000000e+02,1.430000000000000000e+02,1.200000000000000000e+01,8.800000000000000000e+01,1.110000000000000000e+02,1.420000000000000000e+02,7.200000000000000000e+01,6.800000000000000000e+01,8.000000000000000000e+01,1.600000000000000000e+01,1.760000000000000000e+02,1.540000000000000000e+02,7.400000000000000000e+01,6.000000000000000000e+00,1.800000000000000000e+01,1.030000000000000000e+02,7.600000000000000000e+01,4.600000000000000000e+01,2.300000000000000000e+01,3.800000000000000000e+01,7.500000000000000000e+01,9.000000000000000000e+01,1.090000000000000000e+02,1.720000000000000000e+02,8.800000000000000000e+01,1.370000000000000000e+02,1.800000000000000000e+02,2.000000000000000000e+02,2.010000000000000000e+02,1.960000000000000000e+02,1.790000000000000000e+02,1.560000000000000000e+02,1.590000000000000000e+02,1.590000000000000000e+02,1.730000000000000000e+02,1.790000000000000000e+02,1.050000000000000000e+02,1.280000000000000000e+02,1.400000000000000000e+02,1.520000000000000000e+02,1.580000000000000000e+02,1.710000000000000000e+02,1.620000000000000000e+02,1.540000000000000000e+02,1.430000000000000000e+02,1.460000000000000000e+02,1.520000000000000000e+02,1.610000000000000000e+02,1.650000000000000000e+02,1.520000000000000000e+02,1.490000000000000000e+02,1.460000000000000000e+02,1.430000000000000000e+02,1.240000000000000000e+02,1.120000000000000000e+02,8.600000000000000000e+01,6.500000000000000000e+01,5.100000000000000000e+01,4.100000000000000000e+01,5.500000000000000000e+01),
(1.370000000000000000e+02,1.180000000000000000e+02,8.500000000000000000e+01,5.700000000000000000e+01,4.400000000000000000e+01,3.600000000000000000e+01,6.600000000000000000e+01,9.600000000000000000e+01,1.350000000000000000e+02,1.290000000000000000e+02,1.270000000000000000e+02,1.090000000000000000e+02,9.700000000000000000e+01,9.300000000000000000e+01,9.600000000000000000e+01,9.600000000000000000e+01,8.100000000000000000e+01,7.700000000000000000e+01,8.200000000000000000e+01,6.500000000000000000e+01,4.300000000000000000e+01,4.500000000000000000e+01,1.320000000000000000e+02,1.090000000000000000e+02,1.490000000000000000e+02,7.200000000000000000e+01,5.600000000000000000e+01,1.390000000000000000e+02,1.780000000000000000e+02,1.770000000000000000e+02,2.060000000000000000e+02,2.090000000000000000e+02,2.090000000000000000e+02,2.090000000000000000e+02,2.070000000000000000e+02,2.090000000000000000e+02,2.030000000000000000e+02,2.020000000000000000e+02,1.850000000000000000e+02,1.620000000000000000e+02,1.650000000000000000e+02,1.080000000000000000e+02,1.710000000000000000e+02,9.500000000000000000e+01,1.460000000000000000e+02,1.630000000000000000e+02,1.160000000000000000e+02,1.500000000000000000e+02,1.270000000000000000e+02,1.110000000000000000e+02,1.080000000000000000e+02,1.370000000000000000e+02,1.030000000000000000e+02,1.270000000000000000e+02,1.280000000000000000e+02,9.100000000000000000e+01,5.100000000000000000e+01,8.000000000000000000e+01,7.400000000000000000e+01,1.160000000000000000e+02,1.390000000000000000e+02,7.600000000000000000e+01,5.700000000000000000e+01,1.400000000000000000e+01,1.900000000000000000e+01,5.000000000000000000e+00,9.100000000000000000e+01,1.290000000000000000e+02,1.420000000000000000e+02,1.630000000000000000e+02,2.800000000000000000e+01,1.500000000000000000e+01,8.100000000000000000e+01,1.080000000000000000e+02,1.300000000000000000e+02,1.900000000000000000e+01,3.200000000000000000e+01,1.400000000000000000e+01,1.360000000000000000e+02,1.470000000000000000e+02,9.400000000000000000e+01,5.000000000000000000e+00,9.400000000000000000e+01,1.060000000000000000e+02,8.800000000000000000e+01,5.000000000000000000e+01,7.200000000000000000e+01,4.900000000000000000e+01,1.120000000000000000e+02,7.200000000000000000e+01,1.220000000000000000e+02,1.260000000000000000e+02,6.600000000000000000e+01,1.200000000000000000e+02,1.640000000000000000e+02,1.980000000000000000e+02,1.830000000000000000e+02,1.840000000000000000e+02,1.730000000000000000e+02,1.580000000000000000e+02,1.850000000000000000e+02,1.570000000000000000e+02,1.520000000000000000e+02,1.750000000000000000e+02,1.430000000000000000e+02,1.240000000000000000e+02,1.290000000000000000e+02,1.490000000000000000e+02,1.630000000000000000e+02,1.700000000000000000e+02,1.600000000000000000e+02,1.500000000000000000e+02,1.480000000000000000e+02,1.470000000000000000e+02,1.470000000000000000e+02,1.530000000000000000e+02,1.660000000000000000e+02,1.480000000000000000e+02,1.460000000000000000e+02,1.450000000000000000e+02,1.350000000000000000e+02,1.150000000000000000e+02,1.000000000000000000e+02,6.600000000000000000e+01,4.300000000000000000e+01,3.000000000000000000e+01,3.500000000000000000e+01,5.400000000000000000e+01),
(1.370000000000000000e+02,1.210000000000000000e+02,8.600000000000000000e+01,5.900000000000000000e+01,3.400000000000000000e+01,4.200000000000000000e+01,6.700000000000000000e+01,1.010000000000000000e+02,1.320000000000000000e+02,1.230000000000000000e+02,1.180000000000000000e+02,1.030000000000000000e+02,1.030000000000000000e+02,8.700000000000000000e+01,9.600000000000000000e+01,9.600000000000000000e+01,8.400000000000000000e+01,8.600000000000000000e+01,7.800000000000000000e+01,6.900000000000000000e+01,4.300000000000000000e+01,2.200000000000000000e+01,2.200000000000000000e+01,6.900000000000000000e+01,1.160000000000000000e+02,9.100000000000000000e+01,7.000000000000000000e+01,9.600000000000000000e+01,1.650000000000000000e+02,1.920000000000000000e+02,2.090000000000000000e+02,2.090000000000000000e+02,2.090000000000000000e+02,2.060000000000000000e+02,2.010000000000000000e+02,1.960000000000000000e+02,1.930000000000000000e+02,1.860000000000000000e+02,1.800000000000000000e+02,1.940000000000000000e+02,1.530000000000000000e+02,1.570000000000000000e+02,1.570000000000000000e+02,1.250000000000000000e+02,1.010000000000000000e+02,1.650000000000000000e+02,1.190000000000000000e+02,1.590000000000000000e+02,1.390000000000000000e+02,1.200000000000000000e+02,6.200000000000000000e+01,1.050000000000000000e+02,1.030000000000000000e+02,8.100000000000000000e+01,1.110000000000000000e+02,1.160000000000000000e+02,1.260000000000000000e+02,1.280000000000000000e+02,1.610000000000000000e+02,1.300000000000000000e+02,1.530000000000000000e+02,8.100000000000000000e+01,4.700000000000000000e+01,4.000000000000000000e+00,1.200000000000000000e+01,2.000000000000000000e+00,1.070000000000000000e+02,1.270000000000000000e+02,1.380000000000000000e+02,1.760000000000000000e+02,1.300000000000000000e+02,8.000000000000000000e+00,1.400000000000000000e+01,8.100000000000000000e+01,6.800000000000000000e+01,1.200000000000000000e+01,2.000000000000000000e+01,5.000000000000000000e+01,1.000000000000000000e+01,1.080000000000000000e+02,7.800000000000000000e+01,6.000000000000000000e+00,1.400000000000000000e+02,1.760000000000000000e+02,1.090000000000000000e+02,7.900000000000000000e+01,3.800000000000000000e+01,7.200000000000000000e+01,5.900000000000000000e+01,8.000000000000000000e+01,1.270000000000000000e+02,4.900000000000000000e+01,1.100000000000000000e+02,1.230000000000000000e+02,1.790000000000000000e+02,1.730000000000000000e+02,1.560000000000000000e+02,1.730000000000000000e+02,1.570000000000000000e+02,1.680000000000000000e+02,1.580000000000000000e+02,1.360000000000000000e+02,1.460000000000000000e+02,1.760000000000000000e+02,1.760000000000000000e+02,1.250000000000000000e+02,1.350000000000000000e+02,1.470000000000000000e+02,1.620000000000000000e+02,1.680000000000000000e+02,1.590000000000000000e+02,1.450000000000000000e+02,1.420000000000000000e+02,1.400000000000000000e+02,1.480000000000000000e+02,1.540000000000000000e+02,1.590000000000000000e+02,1.510000000000000000e+02,1.480000000000000000e+02,1.460000000000000000e+02,1.330000000000000000e+02,1.150000000000000000e+02,9.700000000000000000e+01,6.900000000000000000e+01,3.800000000000000000e+01,4.100000000000000000e+01,5.400000000000000000e+01,7.300000000000000000e+01),
(1.390000000000000000e+02,1.210000000000000000e+02,8.600000000000000000e+01,5.800000000000000000e+01,3.800000000000000000e+01,3.300000000000000000e+01,6.800000000000000000e+01,9.600000000000000000e+01,1.230000000000000000e+02,1.190000000000000000e+02,1.130000000000000000e+02,1.000000000000000000e+02,9.900000000000000000e+01,9.400000000000000000e+01,9.400000000000000000e+01,1.010000000000000000e+02,8.200000000000000000e+01,7.700000000000000000e+01,7.200000000000000000e+01,7.500000000000000000e+01,5.500000000000000000e+01,4.400000000000000000e+01,4.700000000000000000e+01,3.400000000000000000e+01,8.700000000000000000e+01,8.900000000000000000e+01,6.300000000000000000e+01,8.800000000000000000e+01,1.280000000000000000e+02,1.790000000000000000e+02,1.990000000000000000e+02,2.070000000000000000e+02,2.070000000000000000e+02,2.040000000000000000e+02,2.030000000000000000e+02,1.650000000000000000e+02,1.690000000000000000e+02,1.830000000000000000e+02,1.610000000000000000e+02,1.710000000000000000e+02,1.760000000000000000e+02,1.580000000000000000e+02,1.400000000000000000e+02,1.590000000000000000e+02,1.310000000000000000e+02,1.210000000000000000e+02,1.600000000000000000e+02,1.460000000000000000e+02,1.360000000000000000e+02,1.380000000000000000e+02,8.600000000000000000e+01,6.000000000000000000e+01,6.800000000000000000e+01,1.010000000000000000e+02,8.000000000000000000e+01,1.180000000000000000e+02,1.010000000000000000e+02,1.280000000000000000e+02,1.930000000000000000e+02,1.460000000000000000e+02,1.650000000000000000e+02,1.670000000000000000e+02,6.400000000000000000e+01,6.000000000000000000e+00,6.000000000000000000e+00,4.000000000000000000e+00,5.900000000000000000e+01,1.860000000000000000e+02,1.530000000000000000e+02,1.860000000000000000e+02,1.110000000000000000e+02,1.110000000000000000e+02,1.000000000000000000e+01,1.800000000000000000e+01,3.200000000000000000e+01,2.700000000000000000e+01,6.200000000000000000e+01,2.000000000000000000e+01,8.000000000000000000e+01,5.100000000000000000e+01,5.100000000000000000e+01,5.000000000000000000e+00,9.400000000000000000e+01,1.780000000000000000e+02,1.870000000000000000e+02,8.500000000000000000e+01,1.700000000000000000e+01,1.110000000000000000e+02,7.100000000000000000e+01,1.810000000000000000e+02,7.000000000000000000e+01,7.500000000000000000e+01,1.620000000000000000e+02,1.490000000000000000e+02,1.390000000000000000e+02,1.530000000000000000e+02,1.200000000000000000e+02,1.590000000000000000e+02,1.940000000000000000e+02,1.800000000000000000e+02,1.440000000000000000e+02,1.610000000000000000e+02,1.590000000000000000e+02,1.700000000000000000e+02,1.840000000000000000e+02,1.260000000000000000e+02,1.300000000000000000e+02,1.490000000000000000e+02,1.620000000000000000e+02,1.710000000000000000e+02,1.550000000000000000e+02,1.430000000000000000e+02,1.420000000000000000e+02,1.390000000000000000e+02,1.430000000000000000e+02,1.540000000000000000e+02,1.590000000000000000e+02,1.490000000000000000e+02,1.520000000000000000e+02,1.460000000000000000e+02,1.330000000000000000e+02,1.080000000000000000e+02,9.600000000000000000e+01,6.800000000000000000e+01,4.200000000000000000e+01,5.200000000000000000e+01,7.200000000000000000e+01,9.000000000000000000e+01),
(1.350000000000000000e+02,1.230000000000000000e+02,8.200000000000000000e+01,5.200000000000000000e+01,3.300000000000000000e+01,3.400000000000000000e+01,6.400000000000000000e+01,9.100000000000000000e+01,1.260000000000000000e+02,1.190000000000000000e+02,1.120000000000000000e+02,9.800000000000000000e+01,9.800000000000000000e+01,8.600000000000000000e+01,9.700000000000000000e+01,9.400000000000000000e+01,8.300000000000000000e+01,7.000000000000000000e+01,7.900000000000000000e+01,6.800000000000000000e+01,4.600000000000000000e+01,6.600000000000000000e+01,5.500000000000000000e+01,5.200000000000000000e+01,4.900000000000000000e+01,5.600000000000000000e+01,5.500000000000000000e+01,8.500000000000000000e+01,9.800000000000000000e+01,1.590000000000000000e+02,1.870000000000000000e+02,1.750000000000000000e+02,1.950000000000000000e+02,1.950000000000000000e+02,1.920000000000000000e+02,1.770000000000000000e+02,1.800000000000000000e+02,1.550000000000000000e+02,1.790000000000000000e+02,1.720000000000000000e+02,1.480000000000000000e+02,1.530000000000000000e+02,1.540000000000000000e+02,1.290000000000000000e+02,1.040000000000000000e+02,1.420000000000000000e+02,1.360000000000000000e+02,1.690000000000000000e+02,1.240000000000000000e+02,8.800000000000000000e+01,1.050000000000000000e+02,4.900000000000000000e+01,3.700000000000000000e+01,1.000000000000000000e+01,3.900000000000000000e+01,7.700000000000000000e+01,8.300000000000000000e+01,9.200000000000000000e+01,1.310000000000000000e+02,1.940000000000000000e+02,1.470000000000000000e+02,1.760000000000000000e+02,4.100000000000000000e+01,6.000000000000000000e+00,4.000000000000000000e+00,3.000000000000000000e+00,4.300000000000000000e+01,1.690000000000000000e+02,1.880000000000000000e+02,1.940000000000000000e+02,1.850000000000000000e+02,1.580000000000000000e+02,4.500000000000000000e+01,7.000000000000000000e+00,3.100000000000000000e+01,1.180000000000000000e+02,4.600000000000000000e+01,5.200000000000000000e+01,4.300000000000000000e+01,5.300000000000000000e+01,4.800000000000000000e+01,9.000000000000000000e+00,6.800000000000000000e+01,1.810000000000000000e+02,1.810000000000000000e+02,9.700000000000000000e+01,5.000000000000000000e+00,2.900000000000000000e+01,5.100000000000000000e+01,9.600000000000000000e+01,1.590000000000000000e+02,8.800000000000000000e+01,1.430000000000000000e+02,1.210000000000000000e+02,9.500000000000000000e+01,9.500000000000000000e+01,1.480000000000000000e+02,1.850000000000000000e+02,1.920000000000000000e+02,1.610000000000000000e+02,1.460000000000000000e+02,1.440000000000000000e+02,1.440000000000000000e+02,1.790000000000000000e+02,2.000000000000000000e+02,1.340000000000000000e+02,1.300000000000000000e+02,1.470000000000000000e+02,1.550000000000000000e+02,1.650000000000000000e+02,1.520000000000000000e+02,1.440000000000000000e+02,1.360000000000000000e+02,1.360000000000000000e+02,1.390000000000000000e+02,1.520000000000000000e+02,1.610000000000000000e+02,1.470000000000000000e+02,1.450000000000000000e+02,1.390000000000000000e+02,1.330000000000000000e+02,1.110000000000000000e+02,9.000000000000000000e+01,6.200000000000000000e+01,4.200000000000000000e+01,4.900000000000000000e+01,7.900000000000000000e+01,1.060000000000000000e+02),
(1.330000000000000000e+02,1.190000000000000000e+02,8.200000000000000000e+01,5.700000000000000000e+01,3.600000000000000000e+01,3.200000000000000000e+01,5.800000000000000000e+01,8.700000000000000000e+01,1.130000000000000000e+02,1.160000000000000000e+02,1.100000000000000000e+02,9.900000000000000000e+01,9.400000000000000000e+01,9.000000000000000000e+01,9.200000000000000000e+01,8.900000000000000000e+01,7.600000000000000000e+01,7.800000000000000000e+01,6.400000000000000000e+01,7.700000000000000000e+01,5.700000000000000000e+01,6.400000000000000000e+01,5.600000000000000000e+01,7.500000000000000000e+01,5.000000000000000000e+01,4.900000000000000000e+01,5.400000000000000000e+01,4.900000000000000000e+01,8.200000000000000000e+01,1.510000000000000000e+02,1.950000000000000000e+02,1.990000000000000000e+02,1.680000000000000000e+02,1.100000000000000000e+02,1.460000000000000000e+02,1.710000000000000000e+02,1.520000000000000000e+02,1.850000000000000000e+02,1.950000000000000000e+02,1.390000000000000000e+02,1.400000000000000000e+02,1.400000000000000000e+02,1.140000000000000000e+02,8.900000000000000000e+01,9.200000000000000000e+01,1.280000000000000000e+02,1.090000000000000000e+02,1.480000000000000000e+02,1.290000000000000000e+02,1.150000000000000000e+02,1.410000000000000000e+02,1.300000000000000000e+02,4.900000000000000000e+01,1.000000000000000000e+01,6.000000000000000000e+00,7.000000000000000000e+00,7.000000000000000000e+00,3.900000000000000000e+01,1.170000000000000000e+02,1.770000000000000000e+02,2.100000000000000000e+02,1.600000000000000000e+02,8.700000000000000000e+01,1.300000000000000000e+01,0.000000000000000000e+00,2.000000000000000000e+00,3.400000000000000000e+01,1.970000000000000000e+02,2.000000000000000000e+02,1.990000000000000000e+02,1.720000000000000000e+02,1.570000000000000000e+02,1.370000000000000000e+02,6.600000000000000000e+01,3.300000000000000000e+01,8.200000000000000000e+01,4.200000000000000000e+01,8.800000000000000000e+01,4.500000000000000000e+01,8.500000000000000000e+01,1.100000000000000000e+01,2.700000000000000000e+01,1.100000000000000000e+01,1.190000000000000000e+02,1.850000000000000000e+02,1.490000000000000000e+02,5.500000000000000000e+01,6.000000000000000000e+00,2.400000000000000000e+01,1.230000000000000000e+02,1.340000000000000000e+02,1.640000000000000000e+02,7.600000000000000000e+01,9.500000000000000000e+01,8.300000000000000000e+01,1.210000000000000000e+02,1.380000000000000000e+02,1.350000000000000000e+02,1.500000000000000000e+02,1.210000000000000000e+02,1.500000000000000000e+02,1.520000000000000000e+02,1.370000000000000000e+02,1.930000000000000000e+02,1.820000000000000000e+02,1.090000000000000000e+02,1.260000000000000000e+02,1.470000000000000000e+02,1.540000000000000000e+02,1.640000000000000000e+02,1.500000000000000000e+02,1.420000000000000000e+02,1.340000000000000000e+02,1.350000000000000000e+02,1.440000000000000000e+02,1.530000000000000000e+02,1.540000000000000000e+02,1.480000000000000000e+02,1.430000000000000000e+02,1.390000000000000000e+02,1.320000000000000000e+02,1.030000000000000000e+02,9.200000000000000000e+01,6.700000000000000000e+01,4.300000000000000000e+01,5.200000000000000000e+01,7.600000000000000000e+01,1.040000000000000000e+02),
(1.350000000000000000e+02,1.200000000000000000e+02,8.300000000000000000e+01,5.800000000000000000e+01,3.600000000000000000e+01,2.600000000000000000e+01,5.800000000000000000e+01,8.400000000000000000e+01,1.180000000000000000e+02,1.140000000000000000e+02,1.050000000000000000e+02,9.500000000000000000e+01,8.500000000000000000e+01,9.000000000000000000e+01,8.900000000000000000e+01,9.000000000000000000e+01,8.200000000000000000e+01,7.700000000000000000e+01,7.400000000000000000e+01,7.900000000000000000e+01,7.100000000000000000e+01,7.200000000000000000e+01,9.200000000000000000e+01,1.100000000000000000e+02,6.000000000000000000e+01,6.300000000000000000e+01,4.100000000000000000e+01,5.200000000000000000e+01,9.600000000000000000e+01,1.400000000000000000e+02,1.770000000000000000e+02,1.840000000000000000e+02,1.640000000000000000e+02,1.350000000000000000e+02,1.270000000000000000e+02,1.560000000000000000e+02,1.750000000000000000e+02,1.710000000000000000e+02,1.730000000000000000e+02,1.440000000000000000e+02,1.680000000000000000e+02,1.230000000000000000e+02,8.900000000000000000e+01,1.000000000000000000e+02,1.060000000000000000e+02,1.020000000000000000e+02,1.100000000000000000e+02,1.240000000000000000e+02,1.050000000000000000e+02,1.130000000000000000e+02,1.500000000000000000e+02,1.300000000000000000e+02,8.600000000000000000e+01,1.150000000000000000e+02,5.500000000000000000e+01,5.600000000000000000e+01,1.200000000000000000e+01,1.200000000000000000e+01,8.800000000000000000e+01,1.710000000000000000e+02,1.910000000000000000e+02,2.020000000000000000e+02,1.470000000000000000e+02,1.600000000000000000e+01,1.100000000000000000e+01,3.000000000000000000e+00,1.380000000000000000e+02,1.840000000000000000e+02,1.930000000000000000e+02,1.520000000000000000e+02,1.550000000000000000e+02,1.920000000000000000e+02,1.450000000000000000e+02,1.110000000000000000e+02,1.440000000000000000e+02,7.500000000000000000e+01,5.000000000000000000e+01,8.300000000000000000e+01,1.220000000000000000e+02,1.430000000000000000e+02,7.900000000000000000e+01,2.100000000000000000e+01,2.400000000000000000e+01,1.280000000000000000e+02,1.650000000000000000e+02,1.850000000000000000e+02,1.120000000000000000e+02,7.000000000000000000e+00,6.000000000000000000e+00,9.800000000000000000e+01,1.480000000000000000e+02,8.500000000000000000e+01,9.900000000000000000e+01,4.800000000000000000e+01,9.600000000000000000e+01,1.130000000000000000e+02,1.190000000000000000e+02,1.200000000000000000e+02,1.350000000000000000e+02,1.400000000000000000e+02,1.530000000000000000e+02,1.490000000000000000e+02,1.650000000000000000e+02,1.940000000000000000e+02,1.390000000000000000e+02,9.800000000000000000e+01,1.220000000000000000e+02,1.420000000000000000e+02,1.560000000000000000e+02,1.560000000000000000e+02,1.490000000000000000e+02,1.430000000000000000e+02,1.330000000000000000e+02,1.300000000000000000e+02,1.340000000000000000e+02,1.450000000000000000e+02,1.510000000000000000e+02,1.470000000000000000e+02,1.470000000000000000e+02,1.440000000000000000e+02,1.290000000000000000e+02,1.060000000000000000e+02,8.800000000000000000e+01,6.600000000000000000e+01,4.100000000000000000e+01,4.900000000000000000e+01,7.300000000000000000e+01,1.020000000000000000e+02),
(1.320000000000000000e+02,1.190000000000000000e+02,8.200000000000000000e+01,5.300000000000000000e+01,3.200000000000000000e+01,2.600000000000000000e+01,5.800000000000000000e+01,8.400000000000000000e+01,1.160000000000000000e+02,1.060000000000000000e+02,1.100000000000000000e+02,9.500000000000000000e+01,9.000000000000000000e+01,8.500000000000000000e+01,9.200000000000000000e+01,9.000000000000000000e+01,7.500000000000000000e+01,7.700000000000000000e+01,7.200000000000000000e+01,7.300000000000000000e+01,7.300000000000000000e+01,9.800000000000000000e+01,1.120000000000000000e+02,7.000000000000000000e+01,5.300000000000000000e+01,7.100000000000000000e+01,5.200000000000000000e+01,5.800000000000000000e+01,1.120000000000000000e+02,1.410000000000000000e+02,1.710000000000000000e+02,1.590000000000000000e+02,1.560000000000000000e+02,1.500000000000000000e+02,1.570000000000000000e+02,1.410000000000000000e+02,1.460000000000000000e+02,1.270000000000000000e+02,1.560000000000000000e+02,1.250000000000000000e+02,1.020000000000000000e+02,7.500000000000000000e+01,6.200000000000000000e+01,1.450000000000000000e+02,1.390000000000000000e+02,1.130000000000000000e+02,1.450000000000000000e+02,1.130000000000000000e+02,1.390000000000000000e+02,1.620000000000000000e+02,1.790000000000000000e+02,1.500000000000000000e+02,1.410000000000000000e+02,1.640000000000000000e+02,1.370000000000000000e+02,1.920000000000000000e+02,1.210000000000000000e+02,1.650000000000000000e+02,1.540000000000000000e+02,1.640000000000000000e+02,1.890000000000000000e+02,2.020000000000000000e+02,1.920000000000000000e+02,1.000000000000000000e+02,2.500000000000000000e+01,6.400000000000000000e+01,1.800000000000000000e+02,1.880000000000000000e+02,2.030000000000000000e+02,1.790000000000000000e+02,1.830000000000000000e+02,1.670000000000000000e+02,1.900000000000000000e+02,3.800000000000000000e+01,1.820000000000000000e+02,8.300000000000000000e+01,1.700000000000000000e+02,8.400000000000000000e+01,7.100000000000000000e+01,1.260000000000000000e+02,1.030000000000000000e+02,4.800000000000000000e+01,1.060000000000000000e+02,1.910000000000000000e+02,1.420000000000000000e+02,1.610000000000000000e+02,1.250000000000000000e+02,7.400000000000000000e+01,6.000000000000000000e+00,1.100000000000000000e+01,7.200000000000000000e+01,1.800000000000000000e+02,1.190000000000000000e+02,2.600000000000000000e+01,7.800000000000000000e+01,9.800000000000000000e+01,7.800000000000000000e+01,1.350000000000000000e+02,1.240000000000000000e+02,1.620000000000000000e+02,1.480000000000000000e+02,1.480000000000000000e+02,1.440000000000000000e+02,1.580000000000000000e+02,8.000000000000000000e+01,8.900000000000000000e+01,1.170000000000000000e+02,1.450000000000000000e+02,1.470000000000000000e+02,1.570000000000000000e+02,1.470000000000000000e+02,1.410000000000000000e+02,1.330000000000000000e+02,1.300000000000000000e+02,1.320000000000000000e+02,1.460000000000000000e+02,1.550000000000000000e+02,1.430000000000000000e+02,1.410000000000000000e+02,1.370000000000000000e+02,1.320000000000000000e+02,1.120000000000000000e+02,8.800000000000000000e+01,6.700000000000000000e+01,3.700000000000000000e+01,4.600000000000000000e+01,7.200000000000000000e+01,1.010000000000000000e+02),
(1.290000000000000000e+02,1.130000000000000000e+02,8.400000000000000000e+01,4.500000000000000000e+01,3.200000000000000000e+01,2.900000000000000000e+01,5.800000000000000000e+01,8.200000000000000000e+01,1.170000000000000000e+02,1.070000000000000000e+02,1.080000000000000000e+02,1.000000000000000000e+02,8.900000000000000000e+01,8.300000000000000000e+01,9.300000000000000000e+01,9.600000000000000000e+01,6.900000000000000000e+01,6.800000000000000000e+01,7.900000000000000000e+01,6.700000000000000000e+01,6.700000000000000000e+01,9.700000000000000000e+01,9.200000000000000000e+01,7.900000000000000000e+01,7.100000000000000000e+01,5.200000000000000000e+01,4.600000000000000000e+01,6.800000000000000000e+01,1.130000000000000000e+02,1.510000000000000000e+02,1.540000000000000000e+02,1.660000000000000000e+02,1.550000000000000000e+02,9.300000000000000000e+01,1.340000000000000000e+02,1.780000000000000000e+02,1.380000000000000000e+02,1.660000000000000000e+02,1.110000000000000000e+02,8.200000000000000000e+01,8.600000000000000000e+01,1.030000000000000000e+02,1.240000000000000000e+02,8.300000000000000000e+01,1.480000000000000000e+02,1.110000000000000000e+02,1.580000000000000000e+02,1.640000000000000000e+02,1.650000000000000000e+02,1.990000000000000000e+02,1.970000000000000000e+02,1.890000000000000000e+02,1.690000000000000000e+02,1.910000000000000000e+02,1.700000000000000000e+02,1.970000000000000000e+02,1.640000000000000000e+02,1.680000000000000000e+02,1.870000000000000000e+02,1.970000000000000000e+02,1.700000000000000000e+02,2.070000000000000000e+02,2.020000000000000000e+02,1.940000000000000000e+02,1.410000000000000000e+02,1.140000000000000000e+02,1.760000000000000000e+02,1.760000000000000000e+02,1.880000000000000000e+02,1.870000000000000000e+02,1.860000000000000000e+02,2.060000000000000000e+02,1.620000000000000000e+02,9.200000000000000000e+01,9.500000000000000000e+01,9.700000000000000000e+01,4.500000000000000000e+01,8.900000000000000000e+01,1.070000000000000000e+02,1.670000000000000000e+02,7.300000000000000000e+01,1.150000000000000000e+02,1.090000000000000000e+02,2.000000000000000000e+02,1.600000000000000000e+02,1.570000000000000000e+02,1.640000000000000000e+02,1.660000000000000000e+02,5.000000000000000000e+00,6.000000000000000000e+00,7.300000000000000000e+01,1.890000000000000000e+02,1.350000000000000000e+02,6.100000000000000000e+01,2.800000000000000000e+01,8.000000000000000000e+01,5.000000000000000000e+01,1.040000000000000000e+02,1.250000000000000000e+02,1.520000000000000000e+02,1.330000000000000000e+02,1.480000000000000000e+02,1.660000000000000000e+02,1.160000000000000000e+02,6.700000000000000000e+01,9.100000000000000000e+01,1.170000000000000000e+02,1.390000000000000000e+02,1.490000000000000000e+02,1.540000000000000000e+02,1.470000000000000000e+02,1.410000000000000000e+02,1.310000000000000000e+02,1.260000000000000000e+02,1.390000000000000000e+02,1.420000000000000000e+02,1.570000000000000000e+02,1.470000000000000000e+02,1.430000000000000000e+02,1.410000000000000000e+02,1.260000000000000000e+02,1.100000000000000000e+02,8.900000000000000000e+01,6.400000000000000000e+01,3.900000000000000000e+01,4.500000000000000000e+01,7.000000000000000000e+01,9.600000000000000000e+01),
(1.350000000000000000e+02,1.110000000000000000e+02,7.700000000000000000e+01,4.600000000000000000e+01,2.500000000000000000e+01,2.900000000000000000e+01,5.500000000000000000e+01,8.000000000000000000e+01,1.150000000000000000e+02,1.120000000000000000e+02,1.040000000000000000e+02,1.000000000000000000e+02,8.300000000000000000e+01,7.700000000000000000e+01,7.900000000000000000e+01,8.300000000000000000e+01,6.400000000000000000e+01,5.400000000000000000e+01,7.500000000000000000e+01,7.800000000000000000e+01,6.300000000000000000e+01,7.000000000000000000e+01,8.600000000000000000e+01,7.000000000000000000e+01,7.200000000000000000e+01,7.000000000000000000e+01,6.700000000000000000e+01,1.040000000000000000e+02,1.340000000000000000e+02,1.450000000000000000e+02,1.670000000000000000e+02,1.470000000000000000e+02,1.530000000000000000e+02,1.600000000000000000e+02,1.190000000000000000e+02,1.530000000000000000e+02,1.800000000000000000e+02,1.490000000000000000e+02,7.400000000000000000e+01,9.400000000000000000e+01,1.200000000000000000e+02,8.700000000000000000e+01,1.360000000000000000e+02,1.000000000000000000e+02,1.360000000000000000e+02,1.320000000000000000e+02,1.830000000000000000e+02,1.870000000000000000e+02,1.920000000000000000e+02,2.000000000000000000e+02,2.010000000000000000e+02,1.930000000000000000e+02,2.000000000000000000e+02,1.780000000000000000e+02,1.840000000000000000e+02,1.470000000000000000e+02,1.970000000000000000e+02,1.970000000000000000e+02,1.800000000000000000e+02,2.090000000000000000e+02,2.060000000000000000e+02,2.050000000000000000e+02,2.080000000000000000e+02,2.070000000000000000e+02,2.010000000000000000e+02,2.050000000000000000e+02,2.070000000000000000e+02,1.900000000000000000e+02,1.940000000000000000e+02,1.860000000000000000e+02,1.820000000000000000e+02,1.870000000000000000e+02,1.340000000000000000e+02,1.050000000000000000e+02,1.510000000000000000e+02,1.540000000000000000e+02,9.800000000000000000e+01,1.560000000000000000e+02,6.900000000000000000e+01,1.550000000000000000e+02,9.600000000000000000e+01,4.400000000000000000e+01,1.900000000000000000e+02,1.650000000000000000e+02,1.310000000000000000e+02,1.650000000000000000e+02,1.900000000000000000e+02,2.030000000000000000e+02,5.900000000000000000e+01,1.000000000000000000e+01,1.320000000000000000e+02,1.840000000000000000e+02,1.950000000000000000e+02,4.200000000000000000e+01,9.800000000000000000e+01,1.600000000000000000e+02,1.110000000000000000e+02,9.300000000000000000e+01,1.250000000000000000e+02,1.360000000000000000e+02,1.550000000000000000e+02,1.360000000000000000e+02,9.400000000000000000e+01,5.500000000000000000e+01,6.000000000000000000e+01,9.200000000000000000e+01,1.190000000000000000e+02,1.350000000000000000e+02,1.490000000000000000e+02,1.600000000000000000e+02,1.530000000000000000e+02,1.360000000000000000e+02,1.330000000000000000e+02,1.300000000000000000e+02,1.320000000000000000e+02,1.470000000000000000e+02,1.540000000000000000e+02,1.470000000000000000e+02,1.460000000000000000e+02,1.450000000000000000e+02,1.330000000000000000e+02,1.110000000000000000e+02,8.900000000000000000e+01,6.600000000000000000e+01,4.000000000000000000e+01,4.500000000000000000e+01,7.000000000000000000e+01,9.700000000000000000e+01),
(1.260000000000000000e+02,1.060000000000000000e+02,7.300000000000000000e+01,4.200000000000000000e+01,2.800000000000000000e+01,2.400000000000000000e+01,5.700000000000000000e+01,8.500000000000000000e+01,1.120000000000000000e+02,1.090000000000000000e+02,1.030000000000000000e+02,8.700000000000000000e+01,6.900000000000000000e+01,5.300000000000000000e+01,5.500000000000000000e+01,4.900000000000000000e+01,3.900000000000000000e+01,4.600000000000000000e+01,6.900000000000000000e+01,9.000000000000000000e+01,8.300000000000000000e+01,7.100000000000000000e+01,8.900000000000000000e+01,7.600000000000000000e+01,5.800000000000000000e+01,5.900000000000000000e+01,7.100000000000000000e+01,1.420000000000000000e+02,1.370000000000000000e+02,9.100000000000000000e+01,1.030000000000000000e+02,1.290000000000000000e+02,1.100000000000000000e+02,8.000000000000000000e+01,8.600000000000000000e+01,8.700000000000000000e+01,9.700000000000000000e+01,9.700000000000000000e+01,1.060000000000000000e+02,1.260000000000000000e+02,1.220000000000000000e+02,9.100000000000000000e+01,1.200000000000000000e+02,1.150000000000000000e+02,1.120000000000000000e+02,1.580000000000000000e+02,1.850000000000000000e+02,1.930000000000000000e+02,1.970000000000000000e+02,1.980000000000000000e+02,1.360000000000000000e+02,9.100000000000000000e+01,7.800000000000000000e+01,8.000000000000000000e+00,4.000000000000000000e+00,5.000000000000000000e+00,5.000000000000000000e+00,4.300000000000000000e+01,9.300000000000000000e+01,1.360000000000000000e+02,1.960000000000000000e+02,2.070000000000000000e+02,2.100000000000000000e+02,2.110000000000000000e+02,2.080000000000000000e+02,2.050000000000000000e+02,2.080000000000000000e+02,2.080000000000000000e+02,2.100000000000000000e+02,1.990000000000000000e+02,1.380000000000000000e+02,1.140000000000000000e+02,1.610000000000000000e+02,1.720000000000000000e+02,1.840000000000000000e+02,1.120000000000000000e+02,1.010000000000000000e+02,1.040000000000000000e+02,1.460000000000000000e+02,8.800000000000000000e+01,8.700000000000000000e+01,8.100000000000000000e+01,5.100000000000000000e+01,1.400000000000000000e+02,1.460000000000000000e+02,1.440000000000000000e+02,1.530000000000000000e+02,1.770000000000000000e+02,1.510000000000000000e+02,7.600000000000000000e+01,1.180000000000000000e+02,2.010000000000000000e+02,1.510000000000000000e+02,1.820000000000000000e+02,1.920000000000000000e+02,1.660000000000000000e+02,1.760000000000000000e+02,1.350000000000000000e+02,9.600000000000000000e+01,8.900000000000000000e+01,8.000000000000000000e+01,6.700000000000000000e+01,2.900000000000000000e+01,3.200000000000000000e+01,5.500000000000000000e+01,9.000000000000000000e+01,1.120000000000000000e+02,1.360000000000000000e+02,1.460000000000000000e+02,1.530000000000000000e+02,1.570000000000000000e+02,1.390000000000000000e+02,1.300000000000000000e+02,1.350000000000000000e+02,1.330000000000000000e+02,1.440000000000000000e+02,1.500000000000000000e+02,1.420000000000000000e+02,1.440000000000000000e+02,1.460000000000000000e+02,1.330000000000000000e+02,1.080000000000000000e+02,8.600000000000000000e+01,6.300000000000000000e+01,3.900000000000000000e+01,4.300000000000000000e+01,6.700000000000000000e+01,9.000000000000000000e+01),
(1.290000000000000000e+02,1.100000000000000000e+02,7.200000000000000000e+01,3.900000000000000000e+01,2.300000000000000000e+01,2.700000000000000000e+01,5.400000000000000000e+01,7.900000000000000000e+01,1.050000000000000000e+02,9.500000000000000000e+01,8.900000000000000000e+01,5.900000000000000000e+01,3.600000000000000000e+01,2.700000000000000000e+01,2.800000000000000000e+01,2.900000000000000000e+01,3.700000000000000000e+01,4.700000000000000000e+01,6.500000000000000000e+01,7.600000000000000000e+01,8.700000000000000000e+01,8.300000000000000000e+01,7.400000000000000000e+01,7.800000000000000000e+01,6.600000000000000000e+01,8.200000000000000000e+01,9.300000000000000000e+01,1.560000000000000000e+02,1.310000000000000000e+02,1.000000000000000000e+02,5.100000000000000000e+01,1.220000000000000000e+02,1.470000000000000000e+02,1.310000000000000000e+02,1.100000000000000000e+02,1.670000000000000000e+02,1.560000000000000000e+02,1.170000000000000000e+02,1.420000000000000000e+02,9.900000000000000000e+01,8.400000000000000000e+01,1.090000000000000000e+02,1.050000000000000000e+02,1.250000000000000000e+02,1.420000000000000000e+02,1.390000000000000000e+02,1.500000000000000000e+02,1.550000000000000000e+02,9.100000000000000000e+01,1.600000000000000000e+01,2.000000000000000000e+00,1.000000000000000000e+00,2.000000000000000000e+00,3.000000000000000000e+00,1.000000000000000000e+00,2.000000000000000000e+00,3.000000000000000000e+00,1.000000000000000000e+00,1.000000000000000000e+00,4.000000000000000000e+00,2.000000000000000000e+00,8.500000000000000000e+01,2.040000000000000000e+02,2.090000000000000000e+02,2.120000000000000000e+02,2.100000000000000000e+02,2.110000000000000000e+02,2.110000000000000000e+02,2.100000000000000000e+02,2.050000000000000000e+02,1.380000000000000000e+02,1.840000000000000000e+02,1.850000000000000000e+02,1.820000000000000000e+02,1.300000000000000000e+02,9.000000000000000000e+01,1.740000000000000000e+02,1.340000000000000000e+02,1.580000000000000000e+02,7.900000000000000000e+01,1.080000000000000000e+02,1.740000000000000000e+02,1.410000000000000000e+02,2.300000000000000000e+01,1.430000000000000000e+02,9.000000000000000000e+01,1.690000000000000000e+02,1.740000000000000000e+02,1.970000000000000000e+02,1.870000000000000000e+02,1.900000000000000000e+02,2.070000000000000000e+02,2.050000000000000000e+02,2.060000000000000000e+02,2.080000000000000000e+02,1.880000000000000000e+02,1.680000000000000000e+02,2.030000000000000000e+02,1.870000000000000000e+02,1.500000000000000000e+02,1.140000000000000000e+02,1.050000000000000000e+02,4.500000000000000000e+01,4.400000000000000000e+01,5.300000000000000000e+01,8.200000000000000000e+01,1.070000000000000000e+02,1.350000000000000000e+02,1.430000000000000000e+02,1.560000000000000000e+02,1.490000000000000000e+02,1.410000000000000000e+02,1.350000000000000000e+02,1.350000000000000000e+02,1.290000000000000000e+02,1.430000000000000000e+02,1.450000000000000000e+02,1.350000000000000000e+02,1.370000000000000000e+02,1.390000000000000000e+02,1.320000000000000000e+02,1.100000000000000000e+02,9.100000000000000000e+01,6.500000000000000000e+01,3.800000000000000000e+01,4.300000000000000000e+01,6.700000000000000000e+01,8.900000000000000000e+01),
(1.250000000000000000e+02,9.900000000000000000e+01,7.200000000000000000e+01,4.300000000000000000e+01,2.100000000000000000e+01,2.300000000000000000e+01,4.200000000000000000e+01,6.100000000000000000e+01,8.100000000000000000e+01,7.200000000000000000e+01,5.400000000000000000e+01,3.500000000000000000e+01,1.400000000000000000e+01,1.100000000000000000e+01,1.500000000000000000e+01,1.800000000000000000e+01,1.400000000000000000e+01,3.900000000000000000e+01,7.700000000000000000e+01,6.700000000000000000e+01,6.700000000000000000e+01,5.900000000000000000e+01,8.400000000000000000e+01,7.700000000000000000e+01,6.700000000000000000e+01,9.000000000000000000e+01,1.070000000000000000e+02,1.110000000000000000e+02,1.040000000000000000e+02,9.400000000000000000e+01,7.900000000000000000e+01,5.900000000000000000e+01,1.830000000000000000e+02,1.920000000000000000e+02,9.700000000000000000e+01,1.490000000000000000e+02,1.280000000000000000e+02,1.170000000000000000e+02,6.700000000000000000e+01,8.600000000000000000e+01,1.050000000000000000e+02,9.200000000000000000e+01,1.090000000000000000e+02,1.110000000000000000e+02,1.440000000000000000e+02,1.740000000000000000e+02,1.560000000000000000e+02,8.900000000000000000e+01,2.100000000000000000e+01,7.000000000000000000e+00,2.000000000000000000e+00,6.000000000000000000e+00,9.000000000000000000e+00,1.000000000000000000e+01,8.000000000000000000e+00,9.000000000000000000e+00,6.000000000000000000e+00,2.000000000000000000e+00,2.000000000000000000e+00,2.000000000000000000e+00,3.000000000000000000e+00,5.000000000000000000e+00,5.700000000000000000e+01,1.680000000000000000e+02,2.090000000000000000e+02,2.100000000000000000e+02,2.110000000000000000e+02,2.110000000000000000e+02,2.090000000000000000e+02,2.080000000000000000e+02,1.850000000000000000e+02,1.700000000000000000e+02,1.820000000000000000e+02,1.830000000000000000e+02,8.100000000000000000e+01,1.430000000000000000e+02,1.670000000000000000e+02,1.480000000000000000e+02,1.150000000000000000e+02,1.100000000000000000e+02,1.100000000000000000e+02,7.300000000000000000e+01,1.140000000000000000e+02,8.000000000000000000e+01,1.190000000000000000e+02,1.280000000000000000e+02,1.590000000000000000e+02,1.940000000000000000e+02,2.000000000000000000e+02,2.070000000000000000e+02,2.080000000000000000e+02,2.120000000000000000e+02,2.100000000000000000e+02,2.070000000000000000e+02,1.970000000000000000e+02,1.650000000000000000e+02,1.620000000000000000e+02,1.610000000000000000e+02,1.600000000000000000e+02,1.800000000000000000e+02,1.410000000000000000e+02,6.900000000000000000e+01,3.500000000000000000e+01,3.700000000000000000e+01,5.700000000000000000e+01,8.500000000000000000e+01,1.100000000000000000e+02,1.320000000000000000e+02,1.420000000000000000e+02,1.550000000000000000e+02,1.410000000000000000e+02,1.370000000000000000e+02,1.290000000000000000e+02,1.290000000000000000e+02,1.330000000000000000e+02,1.300000000000000000e+02,1.470000000000000000e+02,1.420000000000000000e+02,1.390000000000000000e+02,1.370000000000000000e+02,1.290000000000000000e+02,1.040000000000000000e+02,8.600000000000000000e+01,6.300000000000000000e+01,3.600000000000000000e+01,3.900000000000000000e+01,6.500000000000000000e+01,8.800000000000000000e+01),
(1.190000000000000000e+02,1.000000000000000000e+02,7.100000000000000000e+01,4.300000000000000000e+01,2.400000000000000000e+01,2.000000000000000000e+01,3.600000000000000000e+01,4.700000000000000000e+01,5.000000000000000000e+01,4.300000000000000000e+01,3.000000000000000000e+01,1.500000000000000000e+01,1.300000000000000000e+01,1.000000000000000000e+01,1.600000000000000000e+01,1.500000000000000000e+01,2.200000000000000000e+01,3.800000000000000000e+01,6.900000000000000000e+01,6.300000000000000000e+01,7.400000000000000000e+01,6.600000000000000000e+01,6.700000000000000000e+01,1.010000000000000000e+02,1.080000000000000000e+02,1.150000000000000000e+02,1.440000000000000000e+02,1.350000000000000000e+02,9.700000000000000000e+01,8.200000000000000000e+01,5.900000000000000000e+01,8.800000000000000000e+01,1.030000000000000000e+02,1.330000000000000000e+02,1.120000000000000000e+02,7.800000000000000000e+01,4.000000000000000000e+01,4.700000000000000000e+01,1.400000000000000000e+01,4.900000000000000000e+01,7.300000000000000000e+01,5.600000000000000000e+01,1.120000000000000000e+02,1.160000000000000000e+02,1.440000000000000000e+02,1.250000000000000000e+02,1.140000000000000000e+02,2.500000000000000000e+01,8.000000000000000000e+00,9.000000000000000000e+00,4.900000000000000000e+01,8.200000000000000000e+01,1.010000000000000000e+02,1.030000000000000000e+02,8.400000000000000000e+01,8.100000000000000000e+01,6.100000000000000000e+01,2.000000000000000000e+01,8.000000000000000000e+00,5.000000000000000000e+00,5.000000000000000000e+00,2.000000000000000000e+00,2.000000000000000000e+00,2.100000000000000000e+01,1.970000000000000000e+02,2.060000000000000000e+02,2.120000000000000000e+02,2.100000000000000000e+02,2.100000000000000000e+02,2.090000000000000000e+02,2.080000000000000000e+02,1.970000000000000000e+02,1.830000000000000000e+02,1.860000000000000000e+02,1.480000000000000000e+02,1.800000000000000000e+02,8.500000000000000000e+01,8.700000000000000000e+01,1.280000000000000000e+02,1.300000000000000000e+02,6.900000000000000000e+01,8.300000000000000000e+01,9.600000000000000000e+01,1.570000000000000000e+02,1.270000000000000000e+02,1.530000000000000000e+02,1.940000000000000000e+02,2.020000000000000000e+02,2.080000000000000000e+02,2.100000000000000000e+02,2.120000000000000000e+02,2.070000000000000000e+02,1.590000000000000000e+02,1.280000000000000000e+02,1.010000000000000000e+02,1.050000000000000000e+02,1.650000000000000000e+02,1.470000000000000000e+02,1.900000000000000000e+02,1.890000000000000000e+02,1.740000000000000000e+02,1.390000000000000000e+02,5.800000000000000000e+01,3.600000000000000000e+01,4.900000000000000000e+01,8.200000000000000000e+01,1.060000000000000000e+02,1.270000000000000000e+02,1.450000000000000000e+02,1.540000000000000000e+02,1.510000000000000000e+02,1.340000000000000000e+02,1.250000000000000000e+02,1.240000000000000000e+02,1.250000000000000000e+02,1.410000000000000000e+02,1.380000000000000000e+02,1.350000000000000000e+02,1.370000000000000000e+02,1.390000000000000000e+02,1.320000000000000000e+02,1.070000000000000000e+02,9.100000000000000000e+01,6.600000000000000000e+01,4.300000000000000000e+01,4.000000000000000000e+01,6.500000000000000000e+01,8.400000000000000000e+01),
(1.190000000000000000e+02,1.060000000000000000e+02,7.100000000000000000e+01,4.000000000000000000e+01,2.600000000000000000e+01,1.800000000000000000e+01,2.500000000000000000e+01,3.800000000000000000e+01,3.400000000000000000e+01,2.300000000000000000e+01,1.700000000000000000e+01,1.400000000000000000e+01,1.500000000000000000e+01,2.300000000000000000e+01,1.800000000000000000e+01,1.600000000000000000e+01,2.800000000000000000e+01,4.700000000000000000e+01,6.200000000000000000e+01,5.800000000000000000e+01,6.500000000000000000e+01,7.700000000000000000e+01,8.800000000000000000e+01,6.500000000000000000e+01,1.210000000000000000e+02,1.260000000000000000e+02,1.470000000000000000e+02,1.240000000000000000e+02,7.800000000000000000e+01,6.200000000000000000e+01,1.000000000000000000e+02,9.500000000000000000e+01,1.290000000000000000e+02,8.600000000000000000e+01,2.100000000000000000e+01,1.700000000000000000e+01,1.000000000000000000e+01,4.000000000000000000e+00,4.000000000000000000e+00,2.000000000000000000e+00,6.000000000000000000e+00,1.300000000000000000e+01,1.400000000000000000e+01,3.800000000000000000e+01,1.260000000000000000e+02,1.750000000000000000e+02,1.780000000000000000e+02,7.600000000000000000e+01,7.000000000000000000e+00,7.800000000000000000e+01,1.390000000000000000e+02,1.750000000000000000e+02,1.580000000000000000e+02,1.460000000000000000e+02,1.610000000000000000e+02,1.740000000000000000e+02,5.800000000000000000e+01,9.700000000000000000e+01,5.100000000000000000e+01,4.100000000000000000e+01,5.300000000000000000e+01,1.000000000000000000e+01,3.000000000000000000e+00,6.000000000000000000e+00,9.900000000000000000e+01,2.100000000000000000e+02,2.100000000000000000e+02,2.120000000000000000e+02,2.110000000000000000e+02,2.100000000000000000e+02,2.090000000000000000e+02,2.010000000000000000e+02,2.010000000000000000e+02,1.840000000000000000e+02,1.830000000000000000e+02,1.590000000000000000e+02,8.500000000000000000e+01,1.590000000000000000e+02,1.070000000000000000e+02,1.190000000000000000e+02,1.240000000000000000e+02,1.150000000000000000e+02,8.900000000000000000e+01,8.000000000000000000e+01,8.400000000000000000e+01,1.270000000000000000e+02,2.060000000000000000e+02,2.050000000000000000e+02,2.020000000000000000e+02,2.050000000000000000e+02,1.500000000000000000e+02,2.500000000000000000e+01,5.000000000000000000e+00,4.000000000000000000e+00,5.000000000000000000e+00,4.000000000000000000e+00,5.000000000000000000e+00,5.000000000000000000e+00,7.000000000000000000e+00,5.800000000000000000e+01,1.080000000000000000e+02,1.360000000000000000e+02,1.000000000000000000e+02,3.800000000000000000e+01,4.400000000000000000e+01,8.100000000000000000e+01,1.060000000000000000e+02,1.300000000000000000e+02,1.360000000000000000e+02,1.450000000000000000e+02,1.450000000000000000e+02,1.270000000000000000e+02,1.230000000000000000e+02,1.240000000000000000e+02,1.280000000000000000e+02,1.350000000000000000e+02,1.440000000000000000e+02,1.320000000000000000e+02,1.350000000000000000e+02,1.360000000000000000e+02,1.240000000000000000e+02,1.050000000000000000e+02,8.600000000000000000e+01,6.400000000000000000e+01,4.100000000000000000e+01,4.400000000000000000e+01,6.800000000000000000e+01,9.000000000000000000e+01),
(1.100000000000000000e+02,8.700000000000000000e+01,5.700000000000000000e+01,3.600000000000000000e+01,2.200000000000000000e+01,1.900000000000000000e+01,2.400000000000000000e+01,2.600000000000000000e+01,2.300000000000000000e+01,1.500000000000000000e+01,1.500000000000000000e+01,1.400000000000000000e+01,2.200000000000000000e+01,2.000000000000000000e+01,1.700000000000000000e+01,1.500000000000000000e+01,1.500000000000000000e+01,4.900000000000000000e+01,7.000000000000000000e+01,7.700000000000000000e+01,6.200000000000000000e+01,6.600000000000000000e+01,1.070000000000000000e+02,8.300000000000000000e+01,9.700000000000000000e+01,1.160000000000000000e+02,1.510000000000000000e+02,8.000000000000000000e+01,5.500000000000000000e+01,6.400000000000000000e+01,7.100000000000000000e+01,7.100000000000000000e+01,7.500000000000000000e+01,2.100000000000000000e+01,1.600000000000000000e+01,6.000000000000000000e+00,5.000000000000000000e+00,3.400000000000000000e+01,3.000000000000000000e+01,6.800000000000000000e+01,3.800000000000000000e+01,4.800000000000000000e+01,1.630000000000000000e+02,1.790000000000000000e+02,1.980000000000000000e+02,1.950000000000000000e+02,1.980000000000000000e+02,1.660000000000000000e+02,1.100000000000000000e+01,1.410000000000000000e+02,1.850000000000000000e+02,2.020000000000000000e+02,2.100000000000000000e+02,1.960000000000000000e+02,1.930000000000000000e+02,2.120000000000000000e+02,1.910000000000000000e+02,1.600000000000000000e+01,1.110000000000000000e+02,8.700000000000000000e+01,1.320000000000000000e+02,1.040000000000000000e+02,2.700000000000000000e+01,5.000000000000000000e+00,1.200000000000000000e+01,1.840000000000000000e+02,2.060000000000000000e+02,2.100000000000000000e+02,2.120000000000000000e+02,2.110000000000000000e+02,2.080000000000000000e+02,1.830000000000000000e+02,1.990000000000000000e+02,1.530000000000000000e+02,1.810000000000000000e+02,1.660000000000000000e+02,1.500000000000000000e+02,1.710000000000000000e+02,1.010000000000000000e+02,1.630000000000000000e+02,7.900000000000000000e+01,4.000000000000000000e+01,7.900000000000000000e+01,9.300000000000000000e+01,8.900000000000000000e+01,1.530000000000000000e+02,2.050000000000000000e+02,2.040000000000000000e+02,1.760000000000000000e+02,4.600000000000000000e+01,2.000000000000000000e+00,0.000000000000000000e+00,2.000000000000000000e+00,4.000000000000000000e+00,5.000000000000000000e+00,5.000000000000000000e+00,5.000000000000000000e+00,2.000000000000000000e+00,4.000000000000000000e+00,2.100000000000000000e+01,8.900000000000000000e+01,1.030000000000000000e+02,5.000000000000000000e+01,5.000000000000000000e+01,5.000000000000000000e+01,9.200000000000000000e+01,9.600000000000000000e+01,1.250000000000000000e+02,1.360000000000000000e+02,1.470000000000000000e+02,1.350000000000000000e+02,1.300000000000000000e+02,1.200000000000000000e+02,1.200000000000000000e+02,1.210000000000000000e+02,1.300000000000000000e+02,1.430000000000000000e+02,1.340000000000000000e+02,1.340000000000000000e+02,1.340000000000000000e+02,1.330000000000000000e+02,1.080000000000000000e+02,8.600000000000000000e+01,6.600000000000000000e+01,4.100000000000000000e+01,4.400000000000000000e+01,6.900000000000000000e+01,8.700000000000000000e+01),
(8.200000000000000000e+01,6.900000000000000000e+01,4.400000000000000000e+01,2.600000000000000000e+01,2.000000000000000000e+01,2.000000000000000000e+01,2.000000000000000000e+01,1.800000000000000000e+01,1.800000000000000000e+01,1.700000000000000000e+01,1.800000000000000000e+01,2.000000000000000000e+01,2.300000000000000000e+01,1.600000000000000000e+01,1.100000000000000000e+01,8.000000000000000000e+00,1.100000000000000000e+01,4.700000000000000000e+01,5.700000000000000000e+01,5.100000000000000000e+01,7.800000000000000000e+01,6.900000000000000000e+01,9.800000000000000000e+01,8.400000000000000000e+01,9.700000000000000000e+01,1.120000000000000000e+02,7.600000000000000000e+01,6.700000000000000000e+01,7.200000000000000000e+01,1.270000000000000000e+02,1.180000000000000000e+02,6.100000000000000000e+01,2.100000000000000000e+01,7.000000000000000000e+00,4.000000000000000000e+00,6.000000000000000000e+00,9.000000000000000000e+00,3.400000000000000000e+01,6.500000000000000000e+01,9.600000000000000000e+01,9.700000000000000000e+01,1.380000000000000000e+02,1.600000000000000000e+02,1.710000000000000000e+02,1.980000000000000000e+02,2.040000000000000000e+02,2.040000000000000000e+02,1.840000000000000000e+02,8.000000000000000000e+00,1.690000000000000000e+02,2.020000000000000000e+02,2.080000000000000000e+02,2.120000000000000000e+02,2.000000000000000000e+02,1.870000000000000000e+02,1.420000000000000000e+02,3.000000000000000000e+00,1.100000000000000000e+01,1.040000000000000000e+02,7.400000000000000000e+01,1.370000000000000000e+02,1.800000000000000000e+02,1.370000000000000000e+02,1.100000000000000000e+01,1.200000000000000000e+01,7.300000000000000000e+01,2.040000000000000000e+02,2.120000000000000000e+02,2.120000000000000000e+02,2.110000000000000000e+02,2.100000000000000000e+02,2.050000000000000000e+02,1.920000000000000000e+02,1.780000000000000000e+02,1.680000000000000000e+02,1.600000000000000000e+02,1.970000000000000000e+02,1.370000000000000000e+02,1.410000000000000000e+02,7.700000000000000000e+01,1.530000000000000000e+02,8.200000000000000000e+01,1.510000000000000000e+02,8.900000000000000000e+01,8.800000000000000000e+01,1.860000000000000000e+02,2.070000000000000000e+02,1.970000000000000000e+02,1.900000000000000000e+01,8.000000000000000000e+00,8.000000000000000000e+00,7.000000000000000000e+00,1.000000000000000000e+01,8.000000000000000000e+00,8.000000000000000000e+00,1.100000000000000000e+01,1.100000000000000000e+01,5.000000000000000000e+00,5.000000000000000000e+00,3.700000000000000000e+01,9.000000000000000000e+01,1.050000000000000000e+02,6.800000000000000000e+01,9.500000000000000000e+01,1.560000000000000000e+02,1.220000000000000000e+02,9.200000000000000000e+01,1.140000000000000000e+02,1.250000000000000000e+02,1.370000000000000000e+02,1.410000000000000000e+02,1.210000000000000000e+02,1.180000000000000000e+02,1.180000000000000000e+02,1.190000000000000000e+02,1.280000000000000000e+02,1.390000000000000000e+02,1.330000000000000000e+02,1.340000000000000000e+02,1.360000000000000000e+02,1.280000000000000000e+02,1.160000000000000000e+02,9.000000000000000000e+01,6.200000000000000000e+01,4.300000000000000000e+01,4.200000000000000000e+01,6.800000000000000000e+01,9.200000000000000000e+01),
(6.000000000000000000e+01,4.600000000000000000e+01,3.500000000000000000e+01,2.700000000000000000e+01,2.000000000000000000e+01,1.600000000000000000e+01,1.400000000000000000e+01,1.300000000000000000e+01,1.300000000000000000e+01,1.600000000000000000e+01,1.800000000000000000e+01,2.400000000000000000e+01,1.700000000000000000e+01,1.300000000000000000e+01,8.000000000000000000e+00,8.000000000000000000e+00,1.300000000000000000e+01,4.200000000000000000e+01,4.600000000000000000e+01,5.800000000000000000e+01,6.300000000000000000e+01,8.300000000000000000e+01,8.200000000000000000e+01,8.200000000000000000e+01,6.900000000000000000e+01,8.700000000000000000e+01,1.160000000000000000e+02,7.100000000000000000e+01,1.060000000000000000e+02,1.210000000000000000e+02,1.440000000000000000e+02,6.200000000000000000e+01,2.500000000000000000e+01,7.000000000000000000e+00,9.000000000000000000e+00,2.900000000000000000e+01,1.900000000000000000e+01,2.200000000000000000e+01,6.300000000000000000e+01,9.100000000000000000e+01,1.150000000000000000e+02,1.280000000000000000e+02,1.420000000000000000e+02,1.840000000000000000e+02,1.950000000000000000e+02,2.070000000000000000e+02,2.090000000000000000e+02,2.060000000000000000e+02,3.900000000000000000e+01,8.000000000000000000e+01,2.040000000000000000e+02,2.120000000000000000e+02,2.040000000000000000e+02,1.970000000000000000e+02,1.880000000000000000e+02,1.380000000000000000e+02,1.000000000000000000e+00,3.700000000000000000e+01,9.000000000000000000e+01,7.900000000000000000e+01,1.290000000000000000e+02,1.810000000000000000e+02,1.970000000000000000e+02,7.500000000000000000e+01,1.300000000000000000e+01,2.800000000000000000e+01,1.850000000000000000e+02,2.130000000000000000e+02,2.120000000000000000e+02,2.120000000000000000e+02,2.100000000000000000e+02,2.000000000000000000e+02,2.010000000000000000e+02,1.910000000000000000e+02,1.810000000000000000e+02,1.870000000000000000e+02,1.130000000000000000e+02,1.600000000000000000e+02,1.820000000000000000e+02,1.250000000000000000e+02,1.380000000000000000e+02,1.000000000000000000e+02,8.100000000000000000e+01,1.480000000000000000e+02,1.140000000000000000e+02,1.820000000000000000e+02,2.120000000000000000e+02,1.530000000000000000e+02,9.000000000000000000e+00,2.130000000000000000e+02,2.150000000000000000e+02,1.430000000000000000e+02,1.700000000000000000e+01,3.500000000000000000e+01,4.400000000000000000e+01,4.100000000000000000e+01,2.400000000000000000e+01,2.300000000000000000e+01,1.000000000000000000e+00,3.700000000000000000e+01,4.900000000000000000e+01,8.700000000000000000e+01,6.600000000000000000e+01,6.100000000000000000e+01,1.500000000000000000e+02,1.160000000000000000e+02,6.500000000000000000e+01,1.040000000000000000e+02,1.260000000000000000e+02,1.380000000000000000e+02,1.320000000000000000e+02,1.200000000000000000e+02,1.180000000000000000e+02,1.130000000000000000e+02,1.120000000000000000e+02,1.270000000000000000e+02,1.360000000000000000e+02,1.290000000000000000e+02,1.350000000000000000e+02,1.330000000000000000e+02,1.270000000000000000e+02,1.110000000000000000e+02,8.500000000000000000e+01,6.200000000000000000e+01,3.800000000000000000e+01,4.600000000000000000e+01,7.100000000000000000e+01,9.200000000000000000e+01),
(2.400000000000000000e+01,2.600000000000000000e+01,2.500000000000000000e+01,2.000000000000000000e+01,1.500000000000000000e+01,1.300000000000000000e+01,1.100000000000000000e+01,1.100000000000000000e+01,1.200000000000000000e+01,1.100000000000000000e+01,1.500000000000000000e+01,2.400000000000000000e+01,1.300000000000000000e+01,9.000000000000000000e+00,1.100000000000000000e+01,1.400000000000000000e+01,1.800000000000000000e+01,4.600000000000000000e+01,3.800000000000000000e+01,4.800000000000000000e+01,6.900000000000000000e+01,6.300000000000000000e+01,5.000000000000000000e+01,4.500000000000000000e+01,3.500000000000000000e+01,5.300000000000000000e+01,1.110000000000000000e+02,1.270000000000000000e+02,1.300000000000000000e+02,1.210000000000000000e+02,9.200000000000000000e+01,1.600000000000000000e+01,1.000000000000000000e+01,1.900000000000000000e+01,1.900000000000000000e+01,1.600000000000000000e+01,2.500000000000000000e+01,7.400000000000000000e+01,9.400000000000000000e+01,6.400000000000000000e+01,9.400000000000000000e+01,6.200000000000000000e+01,1.620000000000000000e+02,1.510000000000000000e+02,1.920000000000000000e+02,2.080000000000000000e+02,2.100000000000000000e+02,2.100000000000000000e+02,1.580000000000000000e+02,7.000000000000000000e+00,1.890000000000000000e+02,2.110000000000000000e+02,2.050000000000000000e+02,1.950000000000000000e+02,1.810000000000000000e+02,1.540000000000000000e+02,6.000000000000000000e+00,1.050000000000000000e+02,7.800000000000000000e+01,9.300000000000000000e+01,1.400000000000000000e+02,1.930000000000000000e+02,2.090000000000000000e+02,5.500000000000000000e+01,1.300000000000000000e+01,1.000000000000000000e+01,5.200000000000000000e+01,2.040000000000000000e+02,2.120000000000000000e+02,2.120000000000000000e+02,2.100000000000000000e+02,2.030000000000000000e+02,1.680000000000000000e+02,1.740000000000000000e+02,1.660000000000000000e+02,1.800000000000000000e+02,1.710000000000000000e+02,1.610000000000000000e+02,1.430000000000000000e+02,1.090000000000000000e+02,1.170000000000000000e+02,1.560000000000000000e+02,1.170000000000000000e+02,1.520000000000000000e+02,7.100000000000000000e+01,2.080000000000000000e+02,2.050000000000000000e+02,5.700000000000000000e+01,1.700000000000000000e+01,2.120000000000000000e+02,1.700000000000000000e+02,2.000000000000000000e+01,1.000000000000000000e+01,5.300000000000000000e+01,4.600000000000000000e+01,6.500000000000000000e+01,7.800000000000000000e+01,4.700000000000000000e+01,1.100000000000000000e+01,1.020000000000000000e+02,1.680000000000000000e+02,1.000000000000000000e+02,4.100000000000000000e+01,1.400000000000000000e+01,2.300000000000000000e+01,5.700000000000000000e+01,6.300000000000000000e+01,9.500000000000000000e+01,1.230000000000000000e+02,1.340000000000000000e+02,1.270000000000000000e+02,1.150000000000000000e+02,1.150000000000000000e+02,1.100000000000000000e+02,1.200000000000000000e+02,1.250000000000000000e+02,1.360000000000000000e+02,1.320000000000000000e+02,1.280000000000000000e+02,1.330000000000000000e+02,1.210000000000000000e+02,1.050000000000000000e+02,8.800000000000000000e+01,6.500000000000000000e+01,4.100000000000000000e+01,4.600000000000000000e+01,6.800000000000000000e+01,9.300000000000000000e+01),
(2.000000000000000000e+01,2.400000000000000000e+01,1.800000000000000000e+01,1.500000000000000000e+01,1.300000000000000000e+01,1.500000000000000000e+01,1.500000000000000000e+01,1.400000000000000000e+01,1.200000000000000000e+01,1.500000000000000000e+01,1.700000000000000000e+01,2.400000000000000000e+01,2.100000000000000000e+01,1.600000000000000000e+01,1.200000000000000000e+01,2.200000000000000000e+01,2.600000000000000000e+01,5.500000000000000000e+01,7.000000000000000000e+01,3.000000000000000000e+01,5.400000000000000000e+01,6.000000000000000000e+01,8.800000000000000000e+01,1.190000000000000000e+02,6.600000000000000000e+01,9.500000000000000000e+01,1.150000000000000000e+02,7.900000000000000000e+01,1.110000000000000000e+02,8.300000000000000000e+01,5.000000000000000000e+01,2.800000000000000000e+01,1.400000000000000000e+01,1.900000000000000000e+01,4.000000000000000000e+01,8.600000000000000000e+01,1.160000000000000000e+02,1.380000000000000000e+02,9.400000000000000000e+01,7.100000000000000000e+01,9.100000000000000000e+01,1.060000000000000000e+02,1.370000000000000000e+02,8.900000000000000000e+01,1.240000000000000000e+02,1.890000000000000000e+02,2.040000000000000000e+02,2.100000000000000000e+02,2.020000000000000000e+02,6.700000000000000000e+01,1.600000000000000000e+01,2.030000000000000000e+02,2.030000000000000000e+02,1.970000000000000000e+02,1.860000000000000000e+02,1.620000000000000000e+02,1.090000000000000000e+02,6.300000000000000000e+01,9.300000000000000000e+01,1.520000000000000000e+02,1.820000000000000000e+02,2.070000000000000000e+02,2.040000000000000000e+02,3.900000000000000000e+01,1.000000000000000000e+01,6.000000000000000000e+00,1.700000000000000000e+01,1.910000000000000000e+02,2.110000000000000000e+02,2.130000000000000000e+02,2.120000000000000000e+02,2.080000000000000000e+02,2.020000000000000000e+02,1.990000000000000000e+02,1.700000000000000000e+02,1.740000000000000000e+02,1.650000000000000000e+02,1.690000000000000000e+02,1.550000000000000000e+02,1.160000000000000000e+02,1.600000000000000000e+02,1.800000000000000000e+02,1.160000000000000000e+02,1.150000000000000000e+02,6.100000000000000000e+01,2.080000000000000000e+02,1.980000000000000000e+02,1.600000000000000000e+01,7.100000000000000000e+01,1.190000000000000000e+02,1.480000000000000000e+02,2.700000000000000000e+01,8.000000000000000000e+00,4.900000000000000000e+01,5.800000000000000000e+01,8.300000000000000000e+01,1.400000000000000000e+02,1.170000000000000000e+02,2.100000000000000000e+01,5.300000000000000000e+01,1.940000000000000000e+02,1.870000000000000000e+02,1.330000000000000000e+02,1.070000000000000000e+02,1.500000000000000000e+01,2.500000000000000000e+01,6.600000000000000000e+01,1.000000000000000000e+02,1.180000000000000000e+02,1.320000000000000000e+02,1.310000000000000000e+02,1.150000000000000000e+02,1.120000000000000000e+02,1.120000000000000000e+02,1.100000000000000000e+02,1.240000000000000000e+02,1.390000000000000000e+02,1.290000000000000000e+02,1.320000000000000000e+02,1.340000000000000000e+02,1.290000000000000000e+02,1.090000000000000000e+02,8.500000000000000000e+01,6.500000000000000000e+01,4.200000000000000000e+01,4.400000000000000000e+01,6.900000000000000000e+01,8.900000000000000000e+01),
(2.400000000000000000e+01,2.900000000000000000e+01,2.100000000000000000e+01,1.500000000000000000e+01,1.000000000000000000e+01,1.500000000000000000e+01,2.000000000000000000e+01,2.300000000000000000e+01,2.000000000000000000e+01,1.800000000000000000e+01,2.500000000000000000e+01,3.000000000000000000e+01,2.600000000000000000e+01,2.600000000000000000e+01,2.100000000000000000e+01,2.500000000000000000e+01,3.300000000000000000e+01,5.100000000000000000e+01,5.100000000000000000e+01,3.400000000000000000e+01,6.700000000000000000e+01,4.200000000000000000e+01,3.700000000000000000e+01,1.000000000000000000e+02,1.000000000000000000e+02,1.100000000000000000e+02,1.110000000000000000e+02,1.340000000000000000e+02,7.800000000000000000e+01,5.400000000000000000e+01,2.200000000000000000e+01,8.000000000000000000e+00,1.800000000000000000e+01,2.900000000000000000e+01,4.800000000000000000e+01,1.370000000000000000e+02,1.710000000000000000e+02,1.550000000000000000e+02,9.900000000000000000e+01,4.900000000000000000e+01,8.800000000000000000e+01,5.500000000000000000e+01,8.900000000000000000e+01,5.600000000000000000e+01,6.300000000000000000e+01,5.800000000000000000e+01,1.710000000000000000e+02,2.060000000000000000e+02,2.050000000000000000e+02,2.020000000000000000e+02,2.700000000000000000e+01,3.700000000000000000e+01,1.710000000000000000e+02,1.910000000000000000e+02,1.840000000000000000e+02,1.840000000000000000e+02,1.260000000000000000e+02,1.190000000000000000e+02,1.520000000000000000e+02,1.870000000000000000e+02,2.020000000000000000e+02,2.080000000000000000e+02,1.200000000000000000e+02,9.000000000000000000e+00,3.000000000000000000e+00,1.600000000000000000e+01,1.300000000000000000e+01,1.320000000000000000e+02,2.050000000000000000e+02,2.120000000000000000e+02,2.140000000000000000e+02,2.090000000000000000e+02,1.650000000000000000e+02,2.070000000000000000e+02,1.960000000000000000e+02,1.840000000000000000e+02,1.800000000000000000e+02,1.600000000000000000e+02,1.360000000000000000e+02,1.470000000000000000e+02,1.360000000000000000e+02,1.220000000000000000e+02,9.200000000000000000e+01,1.380000000000000000e+02,1.110000000000000000e+02,2.060000000000000000e+02,1.810000000000000000e+02,3.300000000000000000e+01,1.280000000000000000e+02,1.690000000000000000e+02,1.810000000000000000e+02,8.600000000000000000e+01,1.600000000000000000e+01,4.700000000000000000e+01,5.600000000000000000e+01,1.230000000000000000e+02,1.550000000000000000e+02,1.630000000000000000e+02,2.600000000000000000e+01,2.300000000000000000e+01,1.890000000000000000e+02,2.010000000000000000e+02,1.860000000000000000e+02,8.100000000000000000e+01,9.000000000000000000e+00,2.200000000000000000e+01,5.600000000000000000e+01,9.500000000000000000e+01,1.100000000000000000e+02,1.290000000000000000e+02,1.260000000000000000e+02,1.170000000000000000e+02,1.080000000000000000e+02,1.080000000000000000e+02,1.110000000000000000e+02,1.260000000000000000e+02,1.350000000000000000e+02,1.300000000000000000e+02,1.330000000000000000e+02,1.330000000000000000e+02,1.290000000000000000e+02,1.090000000000000000e+02,8.800000000000000000e+01,6.500000000000000000e+01,4.300000000000000000e+01,4.600000000000000000e+01,6.700000000000000000e+01,9.300000000000000000e+01),
(2.800000000000000000e+01,2.700000000000000000e+01,1.700000000000000000e+01,8.000000000000000000e+00,1.200000000000000000e+01,1.800000000000000000e+01,2.000000000000000000e+01,2.700000000000000000e+01,3.500000000000000000e+01,3.300000000000000000e+01,3.600000000000000000e+01,3.700000000000000000e+01,3.400000000000000000e+01,3.500000000000000000e+01,3.500000000000000000e+01,2.900000000000000000e+01,3.300000000000000000e+01,4.700000000000000000e+01,4.100000000000000000e+01,5.100000000000000000e+01,5.300000000000000000e+01,4.300000000000000000e+01,2.300000000000000000e+01,8.600000000000000000e+01,9.400000000000000000e+01,6.900000000000000000e+01,9.100000000000000000e+01,4.400000000000000000e+01,5.700000000000000000e+01,2.000000000000000000e+01,1.100000000000000000e+01,9.000000000000000000e+00,4.300000000000000000e+01,1.020000000000000000e+02,9.800000000000000000e+01,1.260000000000000000e+02,1.510000000000000000e+02,1.670000000000000000e+02,1.550000000000000000e+02,1.350000000000000000e+02,1.260000000000000000e+02,6.900000000000000000e+01,3.000000000000000000e+01,4.600000000000000000e+01,4.900000000000000000e+01,1.500000000000000000e+02,7.600000000000000000e+01,1.220000000000000000e+02,1.960000000000000000e+02,2.080000000000000000e+02,1.860000000000000000e+02,2.800000000000000000e+01,8.000000000000000000e+00,8.100000000000000000e+01,1.920000000000000000e+02,2.020000000000000000e+02,1.860000000000000000e+02,1.680000000000000000e+02,2.040000000000000000e+02,1.950000000000000000e+02,1.790000000000000000e+02,1.300000000000000000e+02,3.000000000000000000e+01,2.400000000000000000e+01,1.300000000000000000e+01,6.000000000000000000e+00,6.000000000000000000e+00,4.200000000000000000e+01,1.810000000000000000e+02,2.060000000000000000e+02,2.120000000000000000e+02,2.080000000000000000e+02,1.930000000000000000e+02,2.030000000000000000e+02,1.830000000000000000e+02,2.000000000000000000e+02,1.870000000000000000e+02,2.000000000000000000e+02,1.840000000000000000e+02,1.630000000000000000e+02,1.060000000000000000e+02,1.450000000000000000e+02,1.320000000000000000e+02,1.480000000000000000e+02,5.600000000000000000e+01,1.980000000000000000e+02,1.900000000000000000e+02,4.800000000000000000e+01,1.540000000000000000e+02,1.730000000000000000e+02,1.740000000000000000e+02,1.610000000000000000e+02,7.200000000000000000e+01,3.500000000000000000e+01,7.300000000000000000e+01,1.170000000000000000e+02,1.780000000000000000e+02,1.920000000000000000e+02,9.000000000000000000e+00,3.100000000000000000e+01,1.810000000000000000e+02,2.000000000000000000e+02,1.880000000000000000e+02,9.400000000000000000e+01,2.500000000000000000e+01,2.200000000000000000e+01,5.700000000000000000e+01,9.000000000000000000e+01,1.140000000000000000e+02,1.310000000000000000e+02,1.260000000000000000e+02,1.200000000000000000e+02,1.140000000000000000e+02,1.110000000000000000e+02,1.070000000000000000e+02,1.130000000000000000e+02,1.280000000000000000e+02,1.280000000000000000e+02,1.340000000000000000e+02,1.360000000000000000e+02,1.250000000000000000e+02,1.130000000000000000e+02,9.300000000000000000e+01,6.500000000000000000e+01,4.200000000000000000e+01,4.000000000000000000e+01,6.500000000000000000e+01,8.800000000000000000e+01),
(2.700000000000000000e+01,1.900000000000000000e+01,1.000000000000000000e+01,1.000000000000000000e+01,1.300000000000000000e+01,1.900000000000000000e+01,2.700000000000000000e+01,2.600000000000000000e+01,4.800000000000000000e+01,4.900000000000000000e+01,4.400000000000000000e+01,3.100000000000000000e+01,3.000000000000000000e+01,4.300000000000000000e+01,5.400000000000000000e+01,3.900000000000000000e+01,3.400000000000000000e+01,2.700000000000000000e+01,3.200000000000000000e+01,7.600000000000000000e+01,7.400000000000000000e+01,4.600000000000000000e+01,2.800000000000000000e+01,6.900000000000000000e+01,6.200000000000000000e+01,3.300000000000000000e+01,3.100000000000000000e+01,2.300000000000000000e+01,1.600000000000000000e+01,4.000000000000000000e+00,5.000000000000000000e+00,1.900000000000000000e+01,5.600000000000000000e+01,8.000000000000000000e+01,9.000000000000000000e+01,1.390000000000000000e+02,1.190000000000000000e+02,1.580000000000000000e+02,1.360000000000000000e+02,1.430000000000000000e+02,1.200000000000000000e+02,1.370000000000000000e+02,6.900000000000000000e+01,6.500000000000000000e+01,7.800000000000000000e+01,5.700000000000000000e+01,5.300000000000000000e+01,7.800000000000000000e+01,6.400000000000000000e+01,1.920000000000000000e+02,1.990000000000000000e+02,1.900000000000000000e+02,1.070000000000000000e+02,1.400000000000000000e+01,1.400000000000000000e+01,1.220000000000000000e+02,1.880000000000000000e+02,1.920000000000000000e+02,1.910000000000000000e+02,1.860000000000000000e+02,1.300000000000000000e+02,3.800000000000000000e+01,8.000000000000000000e+00,1.100000000000000000e+01,1.000000000000000000e+01,8.000000000000000000e+00,1.000000000000000000e+01,1.400000000000000000e+01,9.800000000000000000e+01,2.030000000000000000e+02,2.100000000000000000e+02,2.070000000000000000e+02,1.930000000000000000e+02,2.000000000000000000e+02,1.920000000000000000e+02,2.080000000000000000e+02,1.930000000000000000e+02,1.840000000000000000e+02,1.910000000000000000e+02,1.630000000000000000e+02,1.110000000000000000e+02,1.550000000000000000e+02,1.700000000000000000e+02,1.520000000000000000e+02,1.460000000000000000e+02,1.460000000000000000e+02,2.020000000000000000e+02,5.600000000000000000e+01,1.450000000000000000e+02,1.540000000000000000e+02,1.630000000000000000e+02,1.560000000000000000e+02,7.300000000000000000e+01,8.500000000000000000e+01,1.220000000000000000e+02,1.480000000000000000e+02,2.060000000000000000e+02,7.500000000000000000e+01,6.000000000000000000e+00,6.700000000000000000e+01,1.920000000000000000e+02,2.010000000000000000e+02,1.900000000000000000e+02,8.700000000000000000e+01,2.100000000000000000e+01,2.100000000000000000e+01,5.200000000000000000e+01,9.600000000000000000e+01,1.170000000000000000e+02,1.250000000000000000e+02,1.250000000000000000e+02,1.140000000000000000e+02,1.060000000000000000e+02,1.100000000000000000e+02,1.120000000000000000e+02,1.180000000000000000e+02,1.290000000000000000e+02,1.310000000000000000e+02,1.320000000000000000e+02,1.360000000000000000e+02,1.260000000000000000e+02,1.120000000000000000e+02,8.400000000000000000e+01,6.200000000000000000e+01,4.000000000000000000e+01,4.200000000000000000e+01,6.700000000000000000e+01,9.200000000000000000e+01),
(2.200000000000000000e+01,7.000000000000000000e+00,8.000000000000000000e+00,1.500000000000000000e+01,2.500000000000000000e+01,3.200000000000000000e+01,3.800000000000000000e+01,5.000000000000000000e+01,4.700000000000000000e+01,4.800000000000000000e+01,4.300000000000000000e+01,2.800000000000000000e+01,2.900000000000000000e+01,5.300000000000000000e+01,5.500000000000000000e+01,4.200000000000000000e+01,2.800000000000000000e+01,2.600000000000000000e+01,3.700000000000000000e+01,4.700000000000000000e+01,7.200000000000000000e+01,6.000000000000000000e+01,1.800000000000000000e+01,2.000000000000000000e+00,2.500000000000000000e+01,1.500000000000000000e+01,6.000000000000000000e+00,3.000000000000000000e+00,3.000000000000000000e+00,3.000000000000000000e+00,8.000000000000000000e+00,2.400000000000000000e+01,6.900000000000000000e+01,1.380000000000000000e+02,1.430000000000000000e+02,1.440000000000000000e+02,1.530000000000000000e+02,1.530000000000000000e+02,1.120000000000000000e+02,1.720000000000000000e+02,1.490000000000000000e+02,1.440000000000000000e+02,9.700000000000000000e+01,4.300000000000000000e+01,7.300000000000000000e+01,1.780000000000000000e+02,8.800000000000000000e+01,8.900000000000000000e+01,6.200000000000000000e+01,4.000000000000000000e+01,8.900000000000000000e+01,1.790000000000000000e+02,2.090000000000000000e+02,2.020000000000000000e+02,1.080000000000000000e+02,6.600000000000000000e+01,1.100000000000000000e+01,9.000000000000000000e+00,4.000000000000000000e+00,8.000000000000000000e+00,1.100000000000000000e+01,1.400000000000000000e+01,7.700000000000000000e+01,1.030000000000000000e+02,6.900000000000000000e+01,1.800000000000000000e+01,1.800000000000000000e+01,1.400000000000000000e+01,1.700000000000000000e+01,1.220000000000000000e+02,2.050000000000000000e+02,1.880000000000000000e+02,1.640000000000000000e+02,1.860000000000000000e+02,1.950000000000000000e+02,1.930000000000000000e+02,1.840000000000000000e+02,1.820000000000000000e+02,1.970000000000000000e+02,1.660000000000000000e+02,8.400000000000000000e+01,1.360000000000000000e+02,1.410000000000000000e+02,1.330000000000000000e+02,1.680000000000000000e+02,6.300000000000000000e+01,1.890000000000000000e+02,6.100000000000000000e+01,9.800000000000000000e+01,1.420000000000000000e+02,1.490000000000000000e+02,1.790000000000000000e+02,1.220000000000000000e+02,1.410000000000000000e+02,1.660000000000000000e+02,1.790000000000000000e+02,8.200000000000000000e+01,6.000000000000000000e+00,9.000000000000000000e+00,9.700000000000000000e+01,1.810000000000000000e+02,1.990000000000000000e+02,1.420000000000000000e+02,3.100000000000000000e+01,2.600000000000000000e+01,2.400000000000000000e+01,5.600000000000000000e+01,9.400000000000000000e+01,1.050000000000000000e+02,1.220000000000000000e+02,1.220000000000000000e+02,1.130000000000000000e+02,1.050000000000000000e+02,1.060000000000000000e+02,1.060000000000000000e+02,1.220000000000000000e+02,1.290000000000000000e+02,1.270000000000000000e+02,1.390000000000000000e+02,1.320000000000000000e+02,1.260000000000000000e+02,1.100000000000000000e+02,9.100000000000000000e+01,6.500000000000000000e+01,3.900000000000000000e+01,4.300000000000000000e+01,6.500000000000000000e+01,9.300000000000000000e+01),
(1.800000000000000000e+01,9.000000000000000000e+00,1.200000000000000000e+01,2.500000000000000000e+01,4.100000000000000000e+01,5.100000000000000000e+01,5.600000000000000000e+01,5.300000000000000000e+01,4.800000000000000000e+01,3.800000000000000000e+01,3.200000000000000000e+01,2.200000000000000000e+01,1.800000000000000000e+01,2.900000000000000000e+01,3.200000000000000000e+01,2.400000000000000000e+01,3.100000000000000000e+01,6.800000000000000000e+01,6.500000000000000000e+01,9.100000000000000000e+01,6.200000000000000000e+01,3.700000000000000000e+01,3.800000000000000000e+01,1.800000000000000000e+01,4.000000000000000000e+00,5.000000000000000000e+00,3.000000000000000000e+00,4.000000000000000000e+00,4.000000000000000000e+00,6.000000000000000000e+00,1.600000000000000000e+01,2.500000000000000000e+01,6.200000000000000000e+01,1.280000000000000000e+02,1.490000000000000000e+02,1.740000000000000000e+02,1.750000000000000000e+02,1.230000000000000000e+02,1.210000000000000000e+02,1.550000000000000000e+02,1.740000000000000000e+02,1.500000000000000000e+02,1.630000000000000000e+02,5.700000000000000000e+01,8.100000000000000000e+01,8.600000000000000000e+01,1.530000000000000000e+02,8.300000000000000000e+01,1.390000000000000000e+02,7.400000000000000000e+01,7.900000000000000000e+01,8.100000000000000000e+01,6.200000000000000000e+01,1.410000000000000000e+02,1.790000000000000000e+02,1.960000000000000000e+02,2.070000000000000000e+02,1.500000000000000000e+02,1.750000000000000000e+02,1.810000000000000000e+02,1.900000000000000000e+02,2.020000000000000000e+02,2.110000000000000000e+02,2.020000000000000000e+02,1.040000000000000000e+02,6.000000000000000000e+00,1.000000000000000000e+01,5.000000000000000000e+00,2.000000000000000000e+00,1.500000000000000000e+01,7.000000000000000000e+01,1.410000000000000000e+02,1.570000000000000000e+02,1.650000000000000000e+02,1.870000000000000000e+02,1.980000000000000000e+02,1.750000000000000000e+02,1.770000000000000000e+02,1.940000000000000000e+02,1.700000000000000000e+02,1.200000000000000000e+02,1.380000000000000000e+02,1.720000000000000000e+02,1.500000000000000000e+02,1.370000000000000000e+02,6.600000000000000000e+01,9.500000000000000000e+01,4.500000000000000000e+01,5.000000000000000000e+00,3.900000000000000000e+01,1.040000000000000000e+02,1.790000000000000000e+02,1.680000000000000000e+02,1.510000000000000000e+02,8.400000000000000000e+01,2.300000000000000000e+01,9.000000000000000000e+00,1.800000000000000000e+01,7.400000000000000000e+01,1.870000000000000000e+02,1.850000000000000000e+02,1.600000000000000000e+02,5.700000000000000000e+01,3.000000000000000000e+01,5.800000000000000000e+01,3.900000000000000000e+01,7.600000000000000000e+01,1.010000000000000000e+02,1.090000000000000000e+02,1.120000000000000000e+02,1.160000000000000000e+02,1.100000000000000000e+02,1.000000000000000000e+02,1.010000000000000000e+02,1.070000000000000000e+02,1.140000000000000000e+02,1.210000000000000000e+02,1.220000000000000000e+02,1.300000000000000000e+02,1.380000000000000000e+02,1.280000000000000000e+02,1.160000000000000000e+02,9.200000000000000000e+01,6.600000000000000000e+01,4.100000000000000000e+01,3.800000000000000000e+01,5.900000000000000000e+01,8.300000000000000000e+01),
(1.600000000000000000e+01,9.000000000000000000e+00,2.100000000000000000e+01,3.500000000000000000e+01,4.800000000000000000e+01,6.000000000000000000e+01,6.000000000000000000e+01,5.100000000000000000e+01,3.200000000000000000e+01,2.500000000000000000e+01,2.300000000000000000e+01,2.300000000000000000e+01,1.900000000000000000e+01,1.800000000000000000e+01,1.500000000000000000e+01,1.200000000000000000e+01,1.800000000000000000e+01,4.400000000000000000e+01,4.800000000000000000e+01,9.300000000000000000e+01,8.700000000000000000e+01,3.700000000000000000e+01,1.600000000000000000e+01,3.300000000000000000e+01,1.900000000000000000e+01,1.000000000000000000e+01,3.000000000000000000e+00,2.000000000000000000e+00,3.000000000000000000e+00,3.600000000000000000e+01,6.700000000000000000e+01,1.410000000000000000e+02,1.320000000000000000e+02,1.500000000000000000e+02,2.000000000000000000e+02,1.990000000000000000e+02,1.800000000000000000e+02,1.380000000000000000e+02,1.220000000000000000e+02,1.670000000000000000e+02,1.750000000000000000e+02,1.640000000000000000e+02,1.850000000000000000e+02,1.160000000000000000e+02,1.030000000000000000e+02,9.500000000000000000e+01,1.050000000000000000e+02,1.260000000000000000e+02,1.210000000000000000e+02,1.150000000000000000e+02,7.600000000000000000e+01,1.700000000000000000e+02,8.100000000000000000e+01,8.600000000000000000e+01,6.700000000000000000e+01,9.600000000000000000e+01,6.900000000000000000e+01,1.030000000000000000e+02,1.860000000000000000e+02,2.100000000000000000e+02,2.090000000000000000e+02,2.060000000000000000e+02,2.090000000000000000e+02,2.020000000000000000e+02,9.400000000000000000e+01,1.200000000000000000e+01,6.000000000000000000e+00,2.000000000000000000e+00,0.000000000000000000e+00,0.000000000000000000e+00,1.400000000000000000e+01,5.800000000000000000e+01,1.510000000000000000e+02,1.890000000000000000e+02,1.700000000000000000e+02,1.750000000000000000e+02,1.800000000000000000e+02,1.730000000000000000e+02,1.870000000000000000e+02,1.970000000000000000e+02,1.560000000000000000e+02,1.260000000000000000e+02,1.690000000000000000e+02,1.820000000000000000e+02,1.590000000000000000e+02,1.060000000000000000e+02,1.800000000000000000e+01,4.000000000000000000e+00,7.000000000000000000e+00,7.700000000000000000e+01,9.000000000000000000e+01,2.600000000000000000e+01,2.000000000000000000e+01,2.000000000000000000e+01,3.000000000000000000e+01,3.600000000000000000e+01,5.400000000000000000e+01,9.100000000000000000e+01,1.360000000000000000e+02,1.720000000000000000e+02,1.070000000000000000e+02,4.700000000000000000e+01,1.200000000000000000e+01,2.800000000000000000e+01,5.900000000000000000e+01,4.100000000000000000e+01,6.700000000000000000e+01,9.100000000000000000e+01,1.080000000000000000e+02,1.100000000000000000e+02,1.110000000000000000e+02,1.050000000000000000e+02,1.000000000000000000e+02,9.400000000000000000e+01,9.900000000000000000e+01,1.130000000000000000e+02,1.220000000000000000e+02,1.220000000000000000e+02,1.290000000000000000e+02,1.320000000000000000e+02,1.270000000000000000e+02,1.160000000000000000e+02,9.400000000000000000e+01,6.500000000000000000e+01,4.100000000000000000e+01,3.400000000000000000e+01,5.900000000000000000e+01,8.200000000000000000e+01),
(1.500000000000000000e+01,1.300000000000000000e+01,2.300000000000000000e+01,4.500000000000000000e+01,4.800000000000000000e+01,4.800000000000000000e+01,4.400000000000000000e+01,3.300000000000000000e+01,2.400000000000000000e+01,2.400000000000000000e+01,2.500000000000000000e+01,2.500000000000000000e+01,2.100000000000000000e+01,1.400000000000000000e+01,1.200000000000000000e+01,1.300000000000000000e+01,2.400000000000000000e+01,4.000000000000000000e+01,7.500000000000000000e+01,9.700000000000000000e+01,1.210000000000000000e+02,4.700000000000000000e+01,3.300000000000000000e+01,8.900000000000000000e+01,6.400000000000000000e+01,5.900000000000000000e+01,6.000000000000000000e+01,6.300000000000000000e+01,2.800000000000000000e+01,3.700000000000000000e+01,7.700000000000000000e+01,1.250000000000000000e+02,1.490000000000000000e+02,1.810000000000000000e+02,2.000000000000000000e+02,1.970000000000000000e+02,1.780000000000000000e+02,1.440000000000000000e+02,1.470000000000000000e+02,1.160000000000000000e+02,1.370000000000000000e+02,1.550000000000000000e+02,1.120000000000000000e+02,1.820000000000000000e+02,1.710000000000000000e+02,1.520000000000000000e+02,1.030000000000000000e+02,4.500000000000000000e+01,1.430000000000000000e+02,1.800000000000000000e+02,1.110000000000000000e+02,1.420000000000000000e+02,8.900000000000000000e+01,1.480000000000000000e+02,1.710000000000000000e+02,7.300000000000000000e+01,3.900000000000000000e+01,1.020000000000000000e+02,1.200000000000000000e+02,8.300000000000000000e+01,1.630000000000000000e+02,1.530000000000000000e+02,2.000000000000000000e+02,1.890000000000000000e+02,1.510000000000000000e+02,4.100000000000000000e+01,8.000000000000000000e+00,1.200000000000000000e+01,2.000000000000000000e+00,2.000000000000000000e+00,2.000000000000000000e+01,6.100000000000000000e+01,1.260000000000000000e+02,1.540000000000000000e+02,1.460000000000000000e+02,1.560000000000000000e+02,1.690000000000000000e+02,1.840000000000000000e+02,1.810000000000000000e+02,1.760000000000000000e+02,1.740000000000000000e+02,1.660000000000000000e+02,1.460000000000000000e+02,1.910000000000000000e+02,1.720000000000000000e+02,1.380000000000000000e+02,3.200000000000000000e+01,2.000000000000000000e+00,3.000000000000000000e+00,2.500000000000000000e+01,2.000000000000000000e+02,2.030000000000000000e+02,1.970000000000000000e+02,2.030000000000000000e+02,2.060000000000000000e+02,2.020000000000000000e+02,1.570000000000000000e+02,1.630000000000000000e+02,1.650000000000000000e+02,9.800000000000000000e+01,5.500000000000000000e+01,3.100000000000000000e+01,1.700000000000000000e+01,6.200000000000000000e+01,7.400000000000000000e+01,5.100000000000000000e+01,7.100000000000000000e+01,9.000000000000000000e+01,1.050000000000000000e+02,1.060000000000000000e+02,1.140000000000000000e+02,1.030000000000000000e+02,9.100000000000000000e+01,9.300000000000000000e+01,1.000000000000000000e+02,1.120000000000000000e+02,1.180000000000000000e+02,1.210000000000000000e+02,1.230000000000000000e+02,1.320000000000000000e+02,1.250000000000000000e+02,1.120000000000000000e+02,9.400000000000000000e+01,6.800000000000000000e+01,4.100000000000000000e+01,3.900000000000000000e+01,5.900000000000000000e+01,8.100000000000000000e+01),
(1.800000000000000000e+01,2.100000000000000000e+01,3.100000000000000000e+01,4.500000000000000000e+01,4.600000000000000000e+01,3.900000000000000000e+01,2.700000000000000000e+01,2.200000000000000000e+01,1.800000000000000000e+01,2.400000000000000000e+01,2.700000000000000000e+01,2.400000000000000000e+01,1.300000000000000000e+01,1.300000000000000000e+01,1.500000000000000000e+01,1.800000000000000000e+01,2.400000000000000000e+01,3.100000000000000000e+01,8.600000000000000000e+01,9.800000000000000000e+01,6.400000000000000000e+01,6.600000000000000000e+01,2.900000000000000000e+01,9.900000000000000000e+01,1.450000000000000000e+02,1.440000000000000000e+02,9.800000000000000000e+01,1.190000000000000000e+02,7.600000000000000000e+01,1.070000000000000000e+02,1.440000000000000000e+02,1.320000000000000000e+02,1.660000000000000000e+02,1.850000000000000000e+02,1.880000000000000000e+02,1.810000000000000000e+02,2.050000000000000000e+02,1.860000000000000000e+02,1.650000000000000000e+02,1.690000000000000000e+02,1.830000000000000000e+02,1.590000000000000000e+02,1.830000000000000000e+02,1.930000000000000000e+02,1.870000000000000000e+02,1.750000000000000000e+02,1.670000000000000000e+02,1.490000000000000000e+02,1.400000000000000000e+02,1.630000000000000000e+02,1.450000000000000000e+02,1.940000000000000000e+02,1.640000000000000000e+02,1.360000000000000000e+02,1.390000000000000000e+02,1.020000000000000000e+02,1.740000000000000000e+02,1.590000000000000000e+02,1.100000000000000000e+02,8.100000000000000000e+01,1.000000000000000000e+02,9.900000000000000000e+01,1.480000000000000000e+02,1.390000000000000000e+02,1.290000000000000000e+02,1.280000000000000000e+02,4.000000000000000000e+01,1.200000000000000000e+01,8.000000000000000000e+00,1.800000000000000000e+01,5.000000000000000000e+01,1.500000000000000000e+02,1.370000000000000000e+02,1.180000000000000000e+02,1.250000000000000000e+02,1.290000000000000000e+02,1.620000000000000000e+02,1.750000000000000000e+02,1.690000000000000000e+02,1.760000000000000000e+02,1.750000000000000000e+02,1.610000000000000000e+02,1.310000000000000000e+02,1.500000000000000000e+02,1.580000000000000000e+02,1.600000000000000000e+02,1.010000000000000000e+02,1.900000000000000000e+01,0.000000000000000000e+00,1.400000000000000000e+01,1.210000000000000000e+02,2.010000000000000000e+02,1.860000000000000000e+02,1.860000000000000000e+02,1.500000000000000000e+02,9.100000000000000000e+01,7.200000000000000000e+01,9.800000000000000000e+01,9.400000000000000000e+01,3.100000000000000000e+01,2.700000000000000000e+01,1.900000000000000000e+01,3.600000000000000000e+01,7.400000000000000000e+01,4.400000000000000000e+01,3.800000000000000000e+01,6.200000000000000000e+01,8.900000000000000000e+01,9.700000000000000000e+01,1.070000000000000000e+02,1.090000000000000000e+02,9.800000000000000000e+01,9.600000000000000000e+01,9.600000000000000000e+01,1.000000000000000000e+02,1.060000000000000000e+02,1.210000000000000000e+02,1.180000000000000000e+02,1.220000000000000000e+02,1.350000000000000000e+02,1.240000000000000000e+02,1.100000000000000000e+02,9.100000000000000000e+01,7.200000000000000000e+01,4.600000000000000000e+01,3.700000000000000000e+01,5.900000000000000000e+01,8.100000000000000000e+01),
(2.900000000000000000e+01,3.200000000000000000e+01,4.200000000000000000e+01,3.900000000000000000e+01,3.600000000000000000e+01,2.900000000000000000e+01,1.600000000000000000e+01,1.500000000000000000e+01,1.500000000000000000e+01,2.000000000000000000e+01,1.800000000000000000e+01,1.500000000000000000e+01,1.300000000000000000e+01,1.300000000000000000e+01,1.800000000000000000e+01,2.600000000000000000e+01,3.700000000000000000e+01,5.100000000000000000e+01,7.500000000000000000e+01,1.060000000000000000e+02,1.430000000000000000e+02,8.200000000000000000e+01,8.500000000000000000e+01,1.430000000000000000e+02,1.620000000000000000e+02,1.500000000000000000e+02,1.280000000000000000e+02,9.400000000000000000e+01,1.180000000000000000e+02,1.480000000000000000e+02,1.470000000000000000e+02,1.130000000000000000e+02,1.750000000000000000e+02,1.660000000000000000e+02,1.840000000000000000e+02,1.660000000000000000e+02,1.420000000000000000e+02,1.470000000000000000e+02,1.550000000000000000e+02,1.150000000000000000e+02,1.690000000000000000e+02,1.830000000000000000e+02,1.080000000000000000e+02,1.050000000000000000e+02,1.560000000000000000e+02,1.600000000000000000e+02,6.000000000000000000e+01,9.200000000000000000e+01,1.540000000000000000e+02,1.720000000000000000e+02,1.520000000000000000e+02,1.390000000000000000e+02,1.360000000000000000e+02,1.550000000000000000e+02,6.300000000000000000e+01,1.080000000000000000e+02,1.580000000000000000e+02,1.070000000000000000e+02,1.230000000000000000e+02,1.740000000000000000e+02,1.690000000000000000e+02,1.880000000000000000e+02,1.360000000000000000e+02,1.450000000000000000e+02,1.230000000000000000e+02,1.650000000000000000e+02,2.400000000000000000e+01,3.400000000000000000e+01,1.500000000000000000e+01,1.100000000000000000e+01,1.030000000000000000e+02,1.400000000000000000e+02,7.800000000000000000e+01,7.100000000000000000e+01,9.300000000000000000e+01,1.320000000000000000e+02,1.440000000000000000e+02,1.490000000000000000e+02,1.660000000000000000e+02,1.640000000000000000e+02,1.640000000000000000e+02,1.810000000000000000e+02,1.660000000000000000e+02,1.600000000000000000e+02,1.100000000000000000e+02,1.460000000000000000e+02,8.200000000000000000e+01,7.700000000000000000e+01,4.000000000000000000e+00,2.500000000000000000e+01,1.220000000000000000e+02,1.710000000000000000e+02,1.000000000000000000e+02,7.300000000000000000e+01,5.900000000000000000e+01,4.400000000000000000e+01,1.110000000000000000e+02,9.100000000000000000e+01,7.600000000000000000e+01,7.200000000000000000e+01,1.140000000000000000e+02,7.900000000000000000e+01,5.200000000000000000e+01,4.400000000000000000e+01,2.500000000000000000e+01,3.700000000000000000e+01,6.200000000000000000e+01,8.300000000000000000e+01,9.800000000000000000e+01,1.020000000000000000e+02,1.130000000000000000e+02,1.000000000000000000e+02,9.600000000000000000e+01,9.600000000000000000e+01,9.900000000000000000e+01,1.050000000000000000e+02,1.160000000000000000e+02,1.170000000000000000e+02,1.190000000000000000e+02,1.240000000000000000e+02,1.260000000000000000e+02,1.140000000000000000e+02,9.200000000000000000e+01,6.800000000000000000e+01,4.700000000000000000e+01,3.400000000000000000e+01,5.200000000000000000e+01,6.800000000000000000e+01),
(4.700000000000000000e+01,4.600000000000000000e+01,4.100000000000000000e+01,3.900000000000000000e+01,2.500000000000000000e+01,1.500000000000000000e+01,1.500000000000000000e+01,1.600000000000000000e+01,1.900000000000000000e+01,2.000000000000000000e+01,1.600000000000000000e+01,1.300000000000000000e+01,1.900000000000000000e+01,2.400000000000000000e+01,3.400000000000000000e+01,4.200000000000000000e+01,3.800000000000000000e+01,5.700000000000000000e+01,7.800000000000000000e+01,1.280000000000000000e+02,1.600000000000000000e+02,6.900000000000000000e+01,4.700000000000000000e+01,5.700000000000000000e+01,1.390000000000000000e+02,1.810000000000000000e+02,1.670000000000000000e+02,1.380000000000000000e+02,1.470000000000000000e+02,1.680000000000000000e+02,1.720000000000000000e+02,1.760000000000000000e+02,1.640000000000000000e+02,1.660000000000000000e+02,1.670000000000000000e+02,2.000000000000000000e+02,1.910000000000000000e+02,1.580000000000000000e+02,1.800000000000000000e+02,1.810000000000000000e+02,1.940000000000000000e+02,1.870000000000000000e+02,1.420000000000000000e+02,7.700000000000000000e+01,7.300000000000000000e+01,4.400000000000000000e+01,5.100000000000000000e+01,4.900000000000000000e+01,5.700000000000000000e+01,6.000000000000000000e+01,1.190000000000000000e+02,1.600000000000000000e+02,1.580000000000000000e+02,1.220000000000000000e+02,1.380000000000000000e+02,1.230000000000000000e+02,1.450000000000000000e+02,1.490000000000000000e+02,7.800000000000000000e+01,1.320000000000000000e+02,1.760000000000000000e+02,1.150000000000000000e+02,1.630000000000000000e+02,1.310000000000000000e+02,8.800000000000000000e+01,1.450000000000000000e+02,4.800000000000000000e+01,3.400000000000000000e+01,3.700000000000000000e+01,6.300000000000000000e+01,7.900000000000000000e+01,2.300000000000000000e+01,2.200000000000000000e+01,4.700000000000000000e+01,6.000000000000000000e+01,8.200000000000000000e+01,1.160000000000000000e+02,1.530000000000000000e+02,1.550000000000000000e+02,1.710000000000000000e+02,1.740000000000000000e+02,1.690000000000000000e+02,1.740000000000000000e+02,1.650000000000000000e+02,1.730000000000000000e+02,1.370000000000000000e+02,8.600000000000000000e+01,8.200000000000000000e+01,4.600000000000000000e+01,1.900000000000000000e+01,5.700000000000000000e+01,1.330000000000000000e+02,1.070000000000000000e+02,1.670000000000000000e+02,1.070000000000000000e+02,8.300000000000000000e+01,8.900000000000000000e+01,1.000000000000000000e+02,1.710000000000000000e+02,1.200000000000000000e+02,6.000000000000000000e+01,1.070000000000000000e+02,5.100000000000000000e+01,4.300000000000000000e+01,3.300000000000000000e+01,4.900000000000000000e+01,6.800000000000000000e+01,9.200000000000000000e+01,9.900000000000000000e+01,1.170000000000000000e+02,1.210000000000000000e+02,1.070000000000000000e+02,1.020000000000000000e+02,1.010000000000000000e+02,1.000000000000000000e+02,1.080000000000000000e+02,1.190000000000000000e+02,1.170000000000000000e+02,1.190000000000000000e+02,1.240000000000000000e+02,1.230000000000000000e+02,1.090000000000000000e+02,8.900000000000000000e+01,6.400000000000000000e+01,4.200000000000000000e+01,2.500000000000000000e+01,3.800000000000000000e+01,5.300000000000000000e+01),
(4.700000000000000000e+01,4.900000000000000000e+01,2.800000000000000000e+01,1.600000000000000000e+01,1.600000000000000000e+01,1.100000000000000000e+01,1.500000000000000000e+01,2.200000000000000000e+01,2.700000000000000000e+01,2.700000000000000000e+01,2.000000000000000000e+01,2.000000000000000000e+01,3.000000000000000000e+01,4.300000000000000000e+01,4.400000000000000000e+01,6.100000000000000000e+01,6.500000000000000000e+01,7.800000000000000000e+01,1.100000000000000000e+02,1.560000000000000000e+02,1.760000000000000000e+02,1.400000000000000000e+02,5.200000000000000000e+01,2.900000000000000000e+01,9.300000000000000000e+01,1.850000000000000000e+02,2.010000000000000000e+02,1.890000000000000000e+02,1.970000000000000000e+02,1.870000000000000000e+02,1.590000000000000000e+02,1.460000000000000000e+02,1.400000000000000000e+02,1.370000000000000000e+02,1.760000000000000000e+02,1.630000000000000000e+02,1.470000000000000000e+02,1.220000000000000000e+02,1.590000000000000000e+02,1.650000000000000000e+02,1.420000000000000000e+02,1.550000000000000000e+02,1.220000000000000000e+02,1.190000000000000000e+02,1.290000000000000000e+02,1.390000000000000000e+02,8.400000000000000000e+01,1.440000000000000000e+02,1.250000000000000000e+02,1.290000000000000000e+02,1.350000000000000000e+02,1.430000000000000000e+02,1.100000000000000000e+02,9.200000000000000000e+01,6.600000000000000000e+01,1.030000000000000000e+02,1.400000000000000000e+02,1.650000000000000000e+02,1.600000000000000000e+02,1.450000000000000000e+02,1.400000000000000000e+02,1.280000000000000000e+02,1.950000000000000000e+02,1.930000000000000000e+02,1.690000000000000000e+02,9.700000000000000000e+01,9.200000000000000000e+01,1.120000000000000000e+02,6.500000000000000000e+01,1.070000000000000000e+02,2.400000000000000000e+01,1.300000000000000000e+01,4.900000000000000000e+01,3.300000000000000000e+01,3.600000000000000000e+01,6.100000000000000000e+01,1.020000000000000000e+02,1.160000000000000000e+02,1.400000000000000000e+02,1.610000000000000000e+02,1.610000000000000000e+02,1.640000000000000000e+02,1.690000000000000000e+02,1.440000000000000000e+02,1.170000000000000000e+02,1.240000000000000000e+02,8.400000000000000000e+01,4.800000000000000000e+01,5.100000000000000000e+01,3.300000000000000000e+01,7.200000000000000000e+01,9.600000000000000000e+01,1.570000000000000000e+02,1.330000000000000000e+02,1.760000000000000000e+02,1.600000000000000000e+02,1.570000000000000000e+02,5.400000000000000000e+01,8.000000000000000000e+01,7.600000000000000000e+01,7.500000000000000000e+01,8.900000000000000000e+01,3.100000000000000000e+01,5.100000000000000000e+01,2.500000000000000000e+01,3.900000000000000000e+01,6.600000000000000000e+01,8.600000000000000000e+01,1.020000000000000000e+02,1.100000000000000000e+02,1.160000000000000000e+02,1.060000000000000000e+02,1.050000000000000000e+02,1.000000000000000000e+02,1.030000000000000000e+02,1.150000000000000000e+02,1.180000000000000000e+02,1.170000000000000000e+02,1.210000000000000000e+02,1.290000000000000000e+02,1.200000000000000000e+02,1.080000000000000000e+02,8.800000000000000000e+01,6.300000000000000000e+01,3.800000000000000000e+01,2.300000000000000000e+01,2.500000000000000000e+01,3.400000000000000000e+01),
(4.400000000000000000e+01,4.300000000000000000e+01,2.100000000000000000e+01,9.000000000000000000e+00,8.000000000000000000e+00,1.500000000000000000e+01,2.600000000000000000e+01,2.700000000000000000e+01,3.200000000000000000e+01,3.000000000000000000e+01,2.200000000000000000e+01,2.300000000000000000e+01,4.200000000000000000e+01,5.600000000000000000e+01,4.400000000000000000e+01,3.700000000000000000e+01,6.100000000000000000e+01,9.800000000000000000e+01,1.030000000000000000e+02,1.660000000000000000e+02,1.450000000000000000e+02,1.740000000000000000e+02,1.680000000000000000e+02,1.200000000000000000e+02,8.300000000000000000e+01,1.430000000000000000e+02,1.840000000000000000e+02,1.970000000000000000e+02,1.890000000000000000e+02,1.880000000000000000e+02,1.950000000000000000e+02,1.820000000000000000e+02,1.780000000000000000e+02,1.770000000000000000e+02,1.780000000000000000e+02,1.350000000000000000e+02,9.900000000000000000e+01,1.040000000000000000e+02,8.100000000000000000e+01,5.400000000000000000e+01,1.310000000000000000e+02,1.610000000000000000e+02,1.390000000000000000e+02,1.400000000000000000e+02,1.710000000000000000e+02,1.960000000000000000e+02,1.960000000000000000e+02,1.630000000000000000e+02,1.600000000000000000e+02,1.220000000000000000e+02,7.700000000000000000e+01,8.100000000000000000e+01,1.020000000000000000e+02,9.600000000000000000e+01,3.300000000000000000e+01,1.030000000000000000e+02,1.630000000000000000e+02,1.190000000000000000e+02,1.740000000000000000e+02,1.250000000000000000e+02,1.360000000000000000e+02,1.830000000000000000e+02,1.690000000000000000e+02,1.310000000000000000e+02,1.380000000000000000e+02,8.600000000000000000e+01,7.600000000000000000e+01,1.200000000000000000e+02,1.140000000000000000e+02,1.090000000000000000e+02,2.200000000000000000e+01,4.500000000000000000e+01,1.000000000000000000e+01,1.300000000000000000e+01,4.100000000000000000e+01,5.600000000000000000e+01,9.400000000000000000e+01,1.310000000000000000e+02,1.200000000000000000e+02,1.530000000000000000e+02,1.500000000000000000e+02,1.640000000000000000e+02,1.700000000000000000e+02,1.520000000000000000e+02,1.380000000000000000e+02,1.280000000000000000e+02,9.000000000000000000e+01,4.300000000000000000e+01,1.900000000000000000e+01,5.200000000000000000e+01,7.500000000000000000e+01,4.900000000000000000e+01,1.520000000000000000e+02,1.280000000000000000e+02,1.410000000000000000e+02,9.000000000000000000e+01,3.200000000000000000e+01,5.100000000000000000e+01,3.300000000000000000e+01,5.300000000000000000e+01,2.100000000000000000e+01,2.500000000000000000e+01,2.300000000000000000e+01,1.040000000000000000e+02,7.600000000000000000e+01,4.100000000000000000e+01,6.300000000000000000e+01,9.100000000000000000e+01,1.050000000000000000e+02,1.120000000000000000e+02,1.120000000000000000e+02,1.090000000000000000e+02,1.000000000000000000e+02,9.800000000000000000e+01,9.800000000000000000e+01,1.070000000000000000e+02,1.210000000000000000e+02,1.210000000000000000e+02,1.210000000000000000e+02,1.240000000000000000e+02,1.190000000000000000e+02,1.050000000000000000e+02,8.200000000000000000e+01,5.600000000000000000e+01,3.600000000000000000e+01,1.800000000000000000e+01,1.500000000000000000e+01,1.700000000000000000e+01),
(3.900000000000000000e+01,3.100000000000000000e+01,1.800000000000000000e+01,7.000000000000000000e+00,8.000000000000000000e+00,2.100000000000000000e+01,3.400000000000000000e+01,3.300000000000000000e+01,3.000000000000000000e+01,2.400000000000000000e+01,2.300000000000000000e+01,4.200000000000000000e+01,6.600000000000000000e+01,7.200000000000000000e+01,7.500000000000000000e+01,9.500000000000000000e+01,1.140000000000000000e+02,1.280000000000000000e+02,1.450000000000000000e+02,1.500000000000000000e+02,1.330000000000000000e+02,1.850000000000000000e+02,1.370000000000000000e+02,6.500000000000000000e+01,2.100000000000000000e+01,3.600000000000000000e+01,8.800000000000000000e+01,8.800000000000000000e+01,1.560000000000000000e+02,1.660000000000000000e+02,1.410000000000000000e+02,1.360000000000000000e+02,1.750000000000000000e+02,1.570000000000000000e+02,1.290000000000000000e+02,7.400000000000000000e+01,6.800000000000000000e+01,2.300000000000000000e+01,9.000000000000000000e+00,8.000000000000000000e+00,4.000000000000000000e+00,9.000000000000000000e+00,1.700000000000000000e+01,6.400000000000000000e+01,1.080000000000000000e+02,1.210000000000000000e+02,1.500000000000000000e+02,1.350000000000000000e+02,1.240000000000000000e+02,5.700000000000000000e+01,6.500000000000000000e+01,4.700000000000000000e+01,2.600000000000000000e+01,9.900000000000000000e+01,1.080000000000000000e+02,7.200000000000000000e+01,8.100000000000000000e+01,9.400000000000000000e+01,1.010000000000000000e+02,1.230000000000000000e+02,1.510000000000000000e+02,1.790000000000000000e+02,1.860000000000000000e+02,1.740000000000000000e+02,1.440000000000000000e+02,1.830000000000000000e+02,1.320000000000000000e+02,1.110000000000000000e+02,1.070000000000000000e+02,1.180000000000000000e+02,5.200000000000000000e+01,9.000000000000000000e+00,1.300000000000000000e+01,2.900000000000000000e+01,4.400000000000000000e+01,6.700000000000000000e+01,8.900000000000000000e+01,1.190000000000000000e+02,1.010000000000000000e+02,1.120000000000000000e+02,1.500000000000000000e+02,1.370000000000000000e+02,1.440000000000000000e+02,1.780000000000000000e+02,1.540000000000000000e+02,1.210000000000000000e+02,8.900000000000000000e+01,3.900000000000000000e+01,7.000000000000000000e+00,5.400000000000000000e+01,2.800000000000000000e+01,7.800000000000000000e+01,9.700000000000000000e+01,1.300000000000000000e+02,7.100000000000000000e+01,9.200000000000000000e+01,7.600000000000000000e+01,1.090000000000000000e+02,7.300000000000000000e+01,6.300000000000000000e+01,7.600000000000000000e+01,1.400000000000000000e+02,1.270000000000000000e+02,1.080000000000000000e+02,4.800000000000000000e+01,3.600000000000000000e+01,6.300000000000000000e+01,8.700000000000000000e+01,1.050000000000000000e+02,1.150000000000000000e+02,1.150000000000000000e+02,1.090000000000000000e+02,1.050000000000000000e+02,9.900000000000000000e+01,1.010000000000000000e+02,1.070000000000000000e+02,1.150000000000000000e+02,1.170000000000000000e+02,1.170000000000000000e+02,1.140000000000000000e+02,1.110000000000000000e+02,9.800000000000000000e+01,7.600000000000000000e+01,5.400000000000000000e+01,2.700000000000000000e+01,1.200000000000000000e+01,1.000000000000000000e+01,1.000000000000000000e+01),
(3.100000000000000000e+01,2.700000000000000000e+01,2.000000000000000000e+01,1.400000000000000000e+01,1.700000000000000000e+01,3.000000000000000000e+01,4.000000000000000000e+01,3.100000000000000000e+01,2.700000000000000000e+01,3.000000000000000000e+01,3.700000000000000000e+01,6.500000000000000000e+01,7.600000000000000000e+01,6.100000000000000000e+01,4.400000000000000000e+01,3.900000000000000000e+01,5.100000000000000000e+01,6.800000000000000000e+01,1.130000000000000000e+02,1.420000000000000000e+02,1.370000000000000000e+02,1.640000000000000000e+02,1.270000000000000000e+02,7.800000000000000000e+01,3.400000000000000000e+01,1.300000000000000000e+01,1.000000000000000000e+01,3.000000000000000000e+01,3.600000000000000000e+01,4.400000000000000000e+01,2.400000000000000000e+01,6.700000000000000000e+01,6.500000000000000000e+01,5.800000000000000000e+01,3.900000000000000000e+01,1.600000000000000000e+01,1.400000000000000000e+01,9.000000000000000000e+00,5.000000000000000000e+00,5.000000000000000000e+00,1.000000000000000000e+00,4.000000000000000000e+00,1.200000000000000000e+01,6.000000000000000000e+00,9.000000000000000000e+00,1.200000000000000000e+01,2.400000000000000000e+01,7.200000000000000000e+01,7.300000000000000000e+01,3.900000000000000000e+01,7.000000000000000000e+00,6.900000000000000000e+01,3.300000000000000000e+01,3.300000000000000000e+01,9.600000000000000000e+01,1.410000000000000000e+02,1.400000000000000000e+02,1.690000000000000000e+02,1.120000000000000000e+02,1.580000000000000000e+02,1.720000000000000000e+02,1.710000000000000000e+02,1.670000000000000000e+02,1.660000000000000000e+02,1.370000000000000000e+02,1.630000000000000000e+02,1.450000000000000000e+02,1.500000000000000000e+02,1.200000000000000000e+02,1.230000000000000000e+02,7.600000000000000000e+01,3.000000000000000000e+01,3.000000000000000000e+01,1.800000000000000000e+01,6.400000000000000000e+01,6.800000000000000000e+01,8.500000000000000000e+01,8.500000000000000000e+01,8.900000000000000000e+01,9.100000000000000000e+01,1.030000000000000000e+02,9.300000000000000000e+01,1.360000000000000000e+02,1.450000000000000000e+02,1.410000000000000000e+02,1.470000000000000000e+02,1.140000000000000000e+02,6.900000000000000000e+01,9.000000000000000000e+00,5.500000000000000000e+01,6.400000000000000000e+01,9.300000000000000000e+01,1.240000000000000000e+02,1.220000000000000000e+02,1.210000000000000000e+02,1.560000000000000000e+02,7.000000000000000000e+01,8.300000000000000000e+01,6.600000000000000000e+01,4.600000000000000000e+01,8.800000000000000000e+01,1.270000000000000000e+02,1.550000000000000000e+02,9.400000000000000000e+01,5.700000000000000000e+01,4.500000000000000000e+01,6.400000000000000000e+01,9.000000000000000000e+01,9.900000000000000000e+01,1.090000000000000000e+02,1.180000000000000000e+02,1.090000000000000000e+02,1.030000000000000000e+02,9.900000000000000000e+01,1.010000000000000000e+02,1.050000000000000000e+02,1.210000000000000000e+02,1.170000000000000000e+02,1.220000000000000000e+02,1.210000000000000000e+02,1.080000000000000000e+02,8.900000000000000000e+01,7.400000000000000000e+01,4.900000000000000000e+01,2.800000000000000000e+01,1.500000000000000000e+01,1.300000000000000000e+01,1.100000000000000000e+01),
(2.500000000000000000e+01,2.100000000000000000e+01,1.800000000000000000e+01,2.100000000000000000e+01,3.200000000000000000e+01,3.600000000000000000e+01,3.500000000000000000e+01,2.300000000000000000e+01,2.200000000000000000e+01,2.900000000000000000e+01,4.100000000000000000e+01,6.200000000000000000e+01,5.900000000000000000e+01,4.600000000000000000e+01,4.500000000000000000e+01,3.200000000000000000e+01,4.200000000000000000e+01,7.700000000000000000e+01,8.600000000000000000e+01,1.110000000000000000e+02,1.450000000000000000e+02,1.800000000000000000e+02,1.200000000000000000e+02,1.090000000000000000e+02,5.000000000000000000e+01,2.700000000000000000e+01,1.600000000000000000e+01,8.000000000000000000e+00,5.000000000000000000e+00,4.000000000000000000e+00,3.000000000000000000e+00,8.000000000000000000e+00,1.300000000000000000e+01,1.900000000000000000e+01,1.200000000000000000e+01,5.000000000000000000e+00,1.000000000000000000e+01,8.000000000000000000e+00,1.700000000000000000e+01,2.900000000000000000e+01,3.400000000000000000e+01,3.800000000000000000e+01,4.900000000000000000e+01,6.300000000000000000e+01,7.500000000000000000e+01,7.800000000000000000e+01,5.900000000000000000e+01,3.100000000000000000e+01,4.200000000000000000e+01,2.800000000000000000e+01,8.300000000000000000e+01,1.420000000000000000e+02,1.200000000000000000e+02,1.190000000000000000e+02,1.450000000000000000e+02,1.330000000000000000e+02,1.340000000000000000e+02,1.320000000000000000e+02,1.690000000000000000e+02,1.510000000000000000e+02,1.350000000000000000e+02,1.680000000000000000e+02,1.780000000000000000e+02,1.770000000000000000e+02,1.690000000000000000e+02,1.730000000000000000e+02,1.820000000000000000e+02,1.720000000000000000e+02,1.650000000000000000e+02,1.100000000000000000e+02,9.600000000000000000e+01,7.800000000000000000e+01,3.000000000000000000e+01,2.900000000000000000e+01,4.900000000000000000e+01,6.600000000000000000e+01,3.900000000000000000e+01,2.200000000000000000e+01,4.300000000000000000e+01,5.600000000000000000e+01,4.200000000000000000e+01,3.700000000000000000e+01,6.600000000000000000e+01,1.110000000000000000e+02,1.350000000000000000e+02,9.700000000000000000e+01,7.800000000000000000e+01,6.800000000000000000e+01,1.200000000000000000e+01,2.500000000000000000e+01,8.500000000000000000e+01,1.410000000000000000e+02,1.530000000000000000e+02,1.420000000000000000e+02,1.460000000000000000e+02,9.700000000000000000e+01,1.160000000000000000e+02,9.700000000000000000e+01,3.900000000000000000e+01,4.200000000000000000e+01,9.400000000000000000e+01,7.400000000000000000e+01,4.800000000000000000e+01,8.800000000000000000e+01,7.300000000000000000e+01,6.500000000000000000e+01,6.900000000000000000e+01,8.200000000000000000e+01,9.900000000000000000e+01,1.090000000000000000e+02,1.160000000000000000e+02,1.070000000000000000e+02,1.030000000000000000e+02,9.900000000000000000e+01,1.010000000000000000e+02,1.050000000000000000e+02,1.120000000000000000e+02,1.140000000000000000e+02,1.150000000000000000e+02,1.080000000000000000e+02,1.000000000000000000e+02,8.700000000000000000e+01,7.400000000000000000e+01,5.800000000000000000e+01,4.000000000000000000e+01,2.600000000000000000e+01,2.200000000000000000e+01,1.800000000000000000e+01),
(2.300000000000000000e+01,2.800000000000000000e+01,3.000000000000000000e+01,4.100000000000000000e+01,5.300000000000000000e+01,6.100000000000000000e+01,4.800000000000000000e+01,3.500000000000000000e+01,4.100000000000000000e+01,4.600000000000000000e+01,4.900000000000000000e+01,5.100000000000000000e+01,4.900000000000000000e+01,3.300000000000000000e+01,4.700000000000000000e+01,6.400000000000000000e+01,5.200000000000000000e+01,8.900000000000000000e+01,7.900000000000000000e+01,7.800000000000000000e+01,7.500000000000000000e+01,1.760000000000000000e+02,1.650000000000000000e+02,9.900000000000000000e+01,9.800000000000000000e+01,5.600000000000000000e+01,3.800000000000000000e+01,3.400000000000000000e+01,1.500000000000000000e+01,9.000000000000000000e+00,4.000000000000000000e+00,3.000000000000000000e+00,7.000000000000000000e+00,7.000000000000000000e+00,5.000000000000000000e+00,1.700000000000000000e+01,1.300000000000000000e+01,5.000000000000000000e+01,3.100000000000000000e+01,8.600000000000000000e+01,9.600000000000000000e+01,1.320000000000000000e+02,1.410000000000000000e+02,1.400000000000000000e+02,1.530000000000000000e+02,1.150000000000000000e+02,1.140000000000000000e+02,1.010000000000000000e+02,1.010000000000000000e+02,9.900000000000000000e+01,1.130000000000000000e+02,1.530000000000000000e+02,1.720000000000000000e+02,1.290000000000000000e+02,1.250000000000000000e+02,1.570000000000000000e+02,1.420000000000000000e+02,1.320000000000000000e+02,1.170000000000000000e+02,1.660000000000000000e+02,1.520000000000000000e+02,1.540000000000000000e+02,1.580000000000000000e+02,1.510000000000000000e+02,1.940000000000000000e+02,1.970000000000000000e+02,1.600000000000000000e+02,1.800000000000000000e+02,1.770000000000000000e+02,1.730000000000000000e+02,1.650000000000000000e+02,1.370000000000000000e+02,7.900000000000000000e+01,7.000000000000000000e+00,1.800000000000000000e+01,2.100000000000000000e+01,2.000000000000000000e+01,8.100000000000000000e+01,1.240000000000000000e+02,1.130000000000000000e+02,1.160000000000000000e+02,9.500000000000000000e+01,3.800000000000000000e+01,8.500000000000000000e+01,7.300000000000000000e+01,3.200000000000000000e+01,9.000000000000000000e+00,1.400000000000000000e+01,1.300000000000000000e+01,3.900000000000000000e+01,1.100000000000000000e+02,1.330000000000000000e+02,1.330000000000000000e+02,1.230000000000000000e+02,1.560000000000000000e+02,1.160000000000000000e+02,9.700000000000000000e+01,7.800000000000000000e+01,3.400000000000000000e+01,1.600000000000000000e+01,3.600000000000000000e+01,8.000000000000000000e+00,2.300000000000000000e+01,7.700000000000000000e+01,6.700000000000000000e+01,4.800000000000000000e+01,6.700000000000000000e+01,7.800000000000000000e+01,9.800000000000000000e+01,1.080000000000000000e+02,1.130000000000000000e+02,1.090000000000000000e+02,1.010000000000000000e+02,1.000000000000000000e+02,9.600000000000000000e+01,1.050000000000000000e+02,1.110000000000000000e+02,1.130000000000000000e+02,1.060000000000000000e+02,1.020000000000000000e+02,9.000000000000000000e+01,7.700000000000000000e+01,6.900000000000000000e+01,5.400000000000000000e+01,4.200000000000000000e+01,3.100000000000000000e+01,2.600000000000000000e+01,2.700000000000000000e+01),
(3.300000000000000000e+01,4.400000000000000000e+01,5.600000000000000000e+01,7.300000000000000000e+01,8.200000000000000000e+01,7.700000000000000000e+01,7.000000000000000000e+01,6.300000000000000000e+01,7.400000000000000000e+01,7.200000000000000000e+01,6.400000000000000000e+01,6.000000000000000000e+01,3.700000000000000000e+01,3.700000000000000000e+01,7.200000000000000000e+01,8.300000000000000000e+01,6.900000000000000000e+01,8.100000000000000000e+01,9.600000000000000000e+01,9.400000000000000000e+01,6.200000000000000000e+01,1.270000000000000000e+02,1.660000000000000000e+02,1.710000000000000000e+02,1.170000000000000000e+02,8.500000000000000000e+01,3.900000000000000000e+01,2.400000000000000000e+01,8.300000000000000000e+01,5.600000000000000000e+01,7.000000000000000000e+01,6.700000000000000000e+01,3.600000000000000000e+01,2.500000000000000000e+01,2.300000000000000000e+01,4.600000000000000000e+01,8.900000000000000000e+01,8.600000000000000000e+01,1.180000000000000000e+02,1.280000000000000000e+02,1.440000000000000000e+02,1.530000000000000000e+02,1.710000000000000000e+02,1.560000000000000000e+02,9.700000000000000000e+01,2.600000000000000000e+01,5.500000000000000000e+01,7.900000000000000000e+01,1.250000000000000000e+02,1.230000000000000000e+02,1.100000000000000000e+02,1.610000000000000000e+02,1.440000000000000000e+02,1.350000000000000000e+02,1.710000000000000000e+02,1.530000000000000000e+02,1.510000000000000000e+02,1.330000000000000000e+02,1.210000000000000000e+02,1.430000000000000000e+02,8.900000000000000000e+01,1.330000000000000000e+02,1.600000000000000000e+02,1.860000000000000000e+02,1.940000000000000000e+02,1.910000000000000000e+02,1.780000000000000000e+02,1.910000000000000000e+02,1.900000000000000000e+02,2.030000000000000000e+02,2.010000000000000000e+02,2.050000000000000000e+02,1.960000000000000000e+02,3.000000000000000000e+01,2.000000000000000000e+00,1.200000000000000000e+01,9.500000000000000000e+01,1.030000000000000000e+02,1.230000000000000000e+02,1.350000000000000000e+02,1.510000000000000000e+02,1.640000000000000000e+02,1.490000000000000000e+02,1.590000000000000000e+02,1.440000000000000000e+02,1.120000000000000000e+02,6.200000000000000000e+01,2.400000000000000000e+01,9.000000000000000000e+00,7.100000000000000000e+01,8.800000000000000000e+01,1.430000000000000000e+02,1.270000000000000000e+02,1.240000000000000000e+02,1.200000000000000000e+02,1.230000000000000000e+02,1.540000000000000000e+02,4.600000000000000000e+01,1.400000000000000000e+01,5.000000000000000000e+00,2.000000000000000000e+00,3.000000000000000000e+00,1.200000000000000000e+01,4.900000000000000000e+01,5.700000000000000000e+01,4.400000000000000000e+01,6.300000000000000000e+01,8.400000000000000000e+01,1.100000000000000000e+02,1.170000000000000000e+02,1.200000000000000000e+02,1.100000000000000000e+02,1.040000000000000000e+02,1.030000000000000000e+02,1.010000000000000000e+02,1.060000000000000000e+02,1.110000000000000000e+02,1.130000000000000000e+02,1.020000000000000000e+02,9.400000000000000000e+01,8.800000000000000000e+01,7.400000000000000000e+01,6.600000000000000000e+01,6.000000000000000000e+01,5.000000000000000000e+01,4.100000000000000000e+01,4.200000000000000000e+01,3.700000000000000000e+01),
(6.900000000000000000e+01,6.700000000000000000e+01,7.800000000000000000e+01,8.600000000000000000e+01,8.000000000000000000e+01,7.800000000000000000e+01,6.400000000000000000e+01,6.700000000000000000e+01,7.600000000000000000e+01,7.800000000000000000e+01,6.500000000000000000e+01,4.800000000000000000e+01,4.100000000000000000e+01,7.600000000000000000e+01,8.100000000000000000e+01,8.100000000000000000e+01,5.500000000000000000e+01,6.900000000000000000e+01,9.700000000000000000e+01,1.130000000000000000e+02,1.220000000000000000e+02,1.000000000000000000e+02,9.100000000000000000e+01,1.250000000000000000e+02,1.760000000000000000e+02,1.580000000000000000e+02,1.020000000000000000e+02,5.000000000000000000e+01,6.700000000000000000e+01,6.400000000000000000e+01,1.040000000000000000e+02,1.100000000000000000e+02,8.800000000000000000e+01,1.270000000000000000e+02,1.140000000000000000e+02,1.350000000000000000e+02,1.390000000000000000e+02,1.330000000000000000e+02,1.830000000000000000e+02,1.710000000000000000e+02,1.900000000000000000e+02,1.930000000000000000e+02,1.740000000000000000e+02,1.530000000000000000e+02,1.060000000000000000e+02,4.800000000000000000e+01,7.100000000000000000e+01,1.260000000000000000e+02,1.610000000000000000e+02,1.400000000000000000e+02,1.300000000000000000e+02,1.470000000000000000e+02,1.440000000000000000e+02,1.610000000000000000e+02,1.670000000000000000e+02,1.380000000000000000e+02,6.300000000000000000e+01,6.900000000000000000e+01,5.100000000000000000e+01,7.900000000000000000e+01,5.300000000000000000e+01,5.900000000000000000e+01,7.500000000000000000e+01,6.400000000000000000e+01,1.490000000000000000e+02,1.520000000000000000e+02,1.200000000000000000e+02,1.870000000000000000e+02,1.980000000000000000e+02,2.070000000000000000e+02,2.100000000000000000e+02,2.090000000000000000e+02,2.120000000000000000e+02,1.930000000000000000e+02,1.070000000000000000e+02,2.200000000000000000e+01,1.000000000000000000e+01,8.000000000000000000e+00,2.000000000000000000e+00,3.300000000000000000e+01,1.420000000000000000e+02,1.720000000000000000e+02,1.320000000000000000e+02,1.570000000000000000e+02,1.330000000000000000e+02,8.600000000000000000e+01,3.400000000000000000e+01,2.000000000000000000e+01,8.900000000000000000e+01,1.710000000000000000e+02,1.430000000000000000e+02,1.270000000000000000e+02,1.170000000000000000e+02,8.600000000000000000e+01,1.000000000000000000e+02,6.200000000000000000e+01,7.300000000000000000e+01,2.000000000000000000e+01,1.400000000000000000e+01,7.000000000000000000e+00,4.000000000000000000e+00,2.000000000000000000e+00,1.600000000000000000e+01,2.200000000000000000e+01,2.800000000000000000e+01,4.100000000000000000e+01,6.100000000000000000e+01,8.600000000000000000e+01,9.800000000000000000e+01,1.170000000000000000e+02,1.200000000000000000e+02,1.210000000000000000e+02,1.070000000000000000e+02,1.030000000000000000e+02,1.050000000000000000e+02,1.090000000000000000e+02,1.130000000000000000e+02,1.110000000000000000e+02,1.100000000000000000e+02,1.000000000000000000e+02,9.000000000000000000e+01,8.100000000000000000e+01,8.100000000000000000e+01,7.700000000000000000e+01,7.300000000000000000e+01,7.000000000000000000e+01,6.900000000000000000e+01,6.500000000000000000e+01),
(8.000000000000000000e+01,8.500000000000000000e+01,8.400000000000000000e+01,7.700000000000000000e+01,8.100000000000000000e+01,6.600000000000000000e+01,5.600000000000000000e+01,6.200000000000000000e+01,8.400000000000000000e+01,7.900000000000000000e+01,5.500000000000000000e+01,4.000000000000000000e+01,4.800000000000000000e+01,8.300000000000000000e+01,9.300000000000000000e+01,8.700000000000000000e+01,6.900000000000000000e+01,6.900000000000000000e+01,8.700000000000000000e+01,1.290000000000000000e+02,1.060000000000000000e+02,1.190000000000000000e+02,5.900000000000000000e+01,9.400000000000000000e+01,1.730000000000000000e+02,1.680000000000000000e+02,1.020000000000000000e+02,4.500000000000000000e+01,4.000000000000000000e+01,1.510000000000000000e+02,1.780000000000000000e+02,1.270000000000000000e+02,1.210000000000000000e+02,1.740000000000000000e+02,1.820000000000000000e+02,1.580000000000000000e+02,1.450000000000000000e+02,1.620000000000000000e+02,1.740000000000000000e+02,1.950000000000000000e+02,1.770000000000000000e+02,1.790000000000000000e+02,1.750000000000000000e+02,1.650000000000000000e+02,1.620000000000000000e+02,1.580000000000000000e+02,1.520000000000000000e+02,1.430000000000000000e+02,1.530000000000000000e+02,1.630000000000000000e+02,1.320000000000000000e+02,1.450000000000000000e+02,1.860000000000000000e+02,1.760000000000000000e+02,1.670000000000000000e+02,1.370000000000000000e+02,2.800000000000000000e+01,6.400000000000000000e+01,1.400000000000000000e+01,2.500000000000000000e+01,5.500000000000000000e+01,6.000000000000000000e+00,3.000000000000000000e+00,1.800000000000000000e+01,7.600000000000000000e+01,2.600000000000000000e+01,1.000000000000000000e+01,1.320000000000000000e+02,1.710000000000000000e+02,2.090000000000000000e+02,2.110000000000000000e+02,2.110000000000000000e+02,2.120000000000000000e+02,2.100000000000000000e+02,2.110000000000000000e+02,1.720000000000000000e+02,3.400000000000000000e+01,1.200000000000000000e+01,6.000000000000000000e+00,4.000000000000000000e+00,1.150000000000000000e+02,1.440000000000000000e+02,7.900000000000000000e+01,1.360000000000000000e+02,1.030000000000000000e+02,4.000000000000000000e+00,5.000000000000000000e+00,4.500000000000000000e+01,1.970000000000000000e+02,1.950000000000000000e+02,1.270000000000000000e+02,1.010000000000000000e+02,8.400000000000000000e+01,8.300000000000000000e+01,6.100000000000000000e+01,7.600000000000000000e+01,2.700000000000000000e+01,2.600000000000000000e+01,1.300000000000000000e+01,1.100000000000000000e+01,4.000000000000000000e+00,2.000000000000000000e+00,3.000000000000000000e+00,8.000000000000000000e+00,4.000000000000000000e+01,6.700000000000000000e+01,8.400000000000000000e+01,9.700000000000000000e+01,1.070000000000000000e+02,1.200000000000000000e+02,1.180000000000000000e+02,1.130000000000000000e+02,1.120000000000000000e+02,1.070000000000000000e+02,1.100000000000000000e+02,1.080000000000000000e+02,1.130000000000000000e+02,1.150000000000000000e+02,1.110000000000000000e+02,1.010000000000000000e+02,9.400000000000000000e+01,9.500000000000000000e+01,9.300000000000000000e+01,9.100000000000000000e+01,9.400000000000000000e+01,8.800000000000000000e+01,9.000000000000000000e+01,8.500000000000000000e+01),
(8.400000000000000000e+01,9.100000000000000000e+01,8.600000000000000000e+01,7.700000000000000000e+01,7.600000000000000000e+01,5.900000000000000000e+01,5.400000000000000000e+01,7.100000000000000000e+01,6.300000000000000000e+01,5.900000000000000000e+01,4.100000000000000000e+01,4.300000000000000000e+01,7.100000000000000000e+01,1.210000000000000000e+02,9.800000000000000000e+01,9.300000000000000000e+01,8.400000000000000000e+01,7.600000000000000000e+01,7.800000000000000000e+01,6.300000000000000000e+01,1.060000000000000000e+02,1.060000000000000000e+02,1.260000000000000000e+02,1.660000000000000000e+02,1.380000000000000000e+02,1.400000000000000000e+02,9.300000000000000000e+01,9.000000000000000000e+01,5.500000000000000000e+01,8.900000000000000000e+01,1.110000000000000000e+02,1.040000000000000000e+02,1.570000000000000000e+02,1.500000000000000000e+02,1.400000000000000000e+02,1.210000000000000000e+02,1.580000000000000000e+02,1.500000000000000000e+02,9.400000000000000000e+01,1.160000000000000000e+02,1.390000000000000000e+02,1.700000000000000000e+02,1.820000000000000000e+02,1.850000000000000000e+02,1.770000000000000000e+02,1.590000000000000000e+02,1.580000000000000000e+02,1.610000000000000000e+02,1.590000000000000000e+02,1.320000000000000000e+02,1.130000000000000000e+02,9.800000000000000000e+01,8.600000000000000000e+01,1.060000000000000000e+02,1.150000000000000000e+02,1.220000000000000000e+02,1.250000000000000000e+02,1.790000000000000000e+02,5.800000000000000000e+01,9.400000000000000000e+01,1.610000000000000000e+02,1.000000000000000000e+02,2.700000000000000000e+01,1.600000000000000000e+02,1.720000000000000000e+02,6.000000000000000000e+01,9.100000000000000000e+01,1.820000000000000000e+02,2.060000000000000000e+02,2.100000000000000000e+02,2.100000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.100000000000000000e+02,1.830000000000000000e+02,6.900000000000000000e+01,8.000000000000000000e+00,1.300000000000000000e+01,1.170000000000000000e+02,9.600000000000000000e+01,6.100000000000000000e+01,1.070000000000000000e+02,1.200000000000000000e+01,3.200000000000000000e+01,1.630000000000000000e+02,2.090000000000000000e+02,2.080000000000000000e+02,2.040000000000000000e+02,1.670000000000000000e+02,4.100000000000000000e+01,4.800000000000000000e+01,6.000000000000000000e+00,2.000000000000000000e+01,6.200000000000000000e+01,1.900000000000000000e+01,2.000000000000000000e+00,4.000000000000000000e+00,3.000000000000000000e+00,1.000000000000000000e+00,2.000000000000000000e+00,2.000000000000000000e+00,7.000000000000000000e+00,4.500000000000000000e+01,7.100000000000000000e+01,8.200000000000000000e+01,1.020000000000000000e+02,1.190000000000000000e+02,1.230000000000000000e+02,1.190000000000000000e+02,1.120000000000000000e+02,1.040000000000000000e+02,1.010000000000000000e+02,9.800000000000000000e+01,1.060000000000000000e+02,1.160000000000000000e+02,1.180000000000000000e+02,1.150000000000000000e+02,1.060000000000000000e+02,1.010000000000000000e+02,9.600000000000000000e+01,9.600000000000000000e+01,9.600000000000000000e+01,9.700000000000000000e+01,9.900000000000000000e+01,9.500000000000000000e+01,9.600000000000000000e+01),
(7.200000000000000000e+01,9.100000000000000000e+01,7.800000000000000000e+01,7.900000000000000000e+01,6.900000000000000000e+01,5.100000000000000000e+01,4.400000000000000000e+01,4.800000000000000000e+01,4.800000000000000000e+01,3.700000000000000000e+01,3.500000000000000000e+01,7.800000000000000000e+01,1.190000000000000000e+02,1.380000000000000000e+02,1.440000000000000000e+02,1.170000000000000000e+02,7.800000000000000000e+01,1.320000000000000000e+02,1.350000000000000000e+02,8.900000000000000000e+01,9.300000000000000000e+01,1.400000000000000000e+02,1.930000000000000000e+02,1.580000000000000000e+02,1.490000000000000000e+02,1.880000000000000000e+02,1.910000000000000000e+02,1.170000000000000000e+02,8.100000000000000000e+01,7.000000000000000000e+01,9.800000000000000000e+01,1.300000000000000000e+02,1.210000000000000000e+02,1.270000000000000000e+02,1.130000000000000000e+02,1.340000000000000000e+02,7.900000000000000000e+01,7.600000000000000000e+01,8.100000000000000000e+01,8.200000000000000000e+01,1.630000000000000000e+02,2.040000000000000000e+02,2.080000000000000000e+02,2.100000000000000000e+02,2.080000000000000000e+02,2.060000000000000000e+02,1.970000000000000000e+02,1.970000000000000000e+02,1.980000000000000000e+02,2.060000000000000000e+02,2.040000000000000000e+02,2.030000000000000000e+02,2.030000000000000000e+02,2.000000000000000000e+02,1.970000000000000000e+02,1.990000000000000000e+02,1.990000000000000000e+02,2.020000000000000000e+02,1.970000000000000000e+02,2.010000000000000000e+02,2.080000000000000000e+02,2.090000000000000000e+02,1.880000000000000000e+02,1.890000000000000000e+02,1.880000000000000000e+02,1.810000000000000000e+02,1.870000000000000000e+02,2.090000000000000000e+02,2.120000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.110000000000000000e+02,1.500000000000000000e+02,3.900000000000000000e+01,9.800000000000000000e+01,1.170000000000000000e+02,2.700000000000000000e+01,6.500000000000000000e+01,6.300000000000000000e+01,1.100000000000000000e+01,2.050000000000000000e+02,2.100000000000000000e+02,2.140000000000000000e+02,2.110000000000000000e+02,2.010000000000000000e+02,1.610000000000000000e+02,1.400000000000000000e+01,5.300000000000000000e+01,1.300000000000000000e+01,1.100000000000000000e+01,2.300000000000000000e+01,1.200000000000000000e+01,7.000000000000000000e+00,7.000000000000000000e+00,3.000000000000000000e+00,4.000000000000000000e+00,2.000000000000000000e+00,3.000000000000000000e+00,9.000000000000000000e+00,4.600000000000000000e+01,6.100000000000000000e+01,8.400000000000000000e+01,1.050000000000000000e+02,1.100000000000000000e+02,1.120000000000000000e+02,1.060000000000000000e+02,9.900000000000000000e+01,9.900000000000000000e+01,8.800000000000000000e+01,9.200000000000000000e+01,9.700000000000000000e+01,9.900000000000000000e+01,1.120000000000000000e+02,1.070000000000000000e+02,1.050000000000000000e+02,1.040000000000000000e+02,1.000000000000000000e+02,1.040000000000000000e+02,1.010000000000000000e+02,1.000000000000000000e+02,1.060000000000000000e+02,1.030000000000000000e+02,1.030000000000000000e+02),
(8.400000000000000000e+01,8.500000000000000000e+01,7.900000000000000000e+01,7.500000000000000000e+01,7.000000000000000000e+01,4.400000000000000000e+01,3.000000000000000000e+01,3.000000000000000000e+01,4.000000000000000000e+01,4.100000000000000000e+01,3.500000000000000000e+01,7.200000000000000000e+01,1.010000000000000000e+02,1.060000000000000000e+02,1.460000000000000000e+02,1.240000000000000000e+02,7.100000000000000000e+01,7.500000000000000000e+01,1.210000000000000000e+02,1.200000000000000000e+02,1.230000000000000000e+02,1.650000000000000000e+02,1.730000000000000000e+02,1.820000000000000000e+02,1.720000000000000000e+02,1.880000000000000000e+02,1.670000000000000000e+02,1.280000000000000000e+02,1.020000000000000000e+02,9.900000000000000000e+01,1.360000000000000000e+02,1.740000000000000000e+02,2.020000000000000000e+02,1.990000000000000000e+02,1.840000000000000000e+02,1.890000000000000000e+02,1.730000000000000000e+02,1.890000000000000000e+02,1.850000000000000000e+02,1.630000000000000000e+02,1.450000000000000000e+02,1.800000000000000000e+02,1.990000000000000000e+02,2.030000000000000000e+02,2.060000000000000000e+02,2.080000000000000000e+02,2.110000000000000000e+02,2.110000000000000000e+02,2.130000000000000000e+02,2.090000000000000000e+02,2.140000000000000000e+02,2.060000000000000000e+02,2.030000000000000000e+02,1.790000000000000000e+02,1.110000000000000000e+02,9.400000000000000000e+01,1.310000000000000000e+02,1.750000000000000000e+02,1.610000000000000000e+02,1.070000000000000000e+02,1.530000000000000000e+02,1.710000000000000000e+02,8.800000000000000000e+01,8.300000000000000000e+01,1.400000000000000000e+02,1.180000000000000000e+02,6.600000000000000000e+01,1.540000000000000000e+02,1.880000000000000000e+02,1.940000000000000000e+02,2.110000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.120000000000000000e+02,2.070000000000000000e+02,1.400000000000000000e+01,3.600000000000000000e+01,5.100000000000000000e+01,3.000000000000000000e+00,3.200000000000000000e+01,1.800000000000000000e+01,1.180000000000000000e+02,2.130000000000000000e+02,2.120000000000000000e+02,2.120000000000000000e+02,2.100000000000000000e+02,2.010000000000000000e+02,1.690000000000000000e+02,1.140000000000000000e+02,1.180000000000000000e+02,1.310000000000000000e+02,7.100000000000000000e+01,3.800000000000000000e+01,1.500000000000000000e+01,1.400000000000000000e+01,1.700000000000000000e+01,1.700000000000000000e+01,2.100000000000000000e+01,1.300000000000000000e+01,1.100000000000000000e+01,1.600000000000000000e+01,4.900000000000000000e+01,7.100000000000000000e+01,7.800000000000000000e+01,9.000000000000000000e+01,9.100000000000000000e+01,8.900000000000000000e+01,8.800000000000000000e+01,8.100000000000000000e+01,7.200000000000000000e+01,7.300000000000000000e+01,7.500000000000000000e+01,7.500000000000000000e+01,8.100000000000000000e+01,8.700000000000000000e+01,8.900000000000000000e+01,9.100000000000000000e+01,8.500000000000000000e+01,8.900000000000000000e+01,9.000000000000000000e+01,9.000000000000000000e+01,9.100000000000000000e+01,9.100000000000000000e+01,9.200000000000000000e+01,9.000000000000000000e+01),
(8.500000000000000000e+01,7.500000000000000000e+01,7.000000000000000000e+01,6.900000000000000000e+01,5.900000000000000000e+01,4.000000000000000000e+01,2.900000000000000000e+01,2.300000000000000000e+01,5.900000000000000000e+01,9.300000000000000000e+01,7.200000000000000000e+01,6.800000000000000000e+01,7.300000000000000000e+01,9.600000000000000000e+01,1.110000000000000000e+02,1.410000000000000000e+02,1.300000000000000000e+02,8.800000000000000000e+01,6.300000000000000000e+01,7.600000000000000000e+01,6.700000000000000000e+01,8.200000000000000000e+01,1.300000000000000000e+02,1.780000000000000000e+02,1.770000000000000000e+02,1.960000000000000000e+02,1.950000000000000000e+02,1.770000000000000000e+02,1.150000000000000000e+02,7.800000000000000000e+01,4.500000000000000000e+01,2.500000000000000000e+01,6.900000000000000000e+01,9.600000000000000000e+01,1.200000000000000000e+02,1.130000000000000000e+02,6.700000000000000000e+01,4.800000000000000000e+01,8.000000000000000000e+01,1.260000000000000000e+02,1.610000000000000000e+02,1.900000000000000000e+02,1.990000000000000000e+02,2.030000000000000000e+02,2.050000000000000000e+02,1.970000000000000000e+02,1.610000000000000000e+02,1.510000000000000000e+02,1.510000000000000000e+02,1.710000000000000000e+02,1.770000000000000000e+02,1.690000000000000000e+02,1.400000000000000000e+02,1.410000000000000000e+02,1.870000000000000000e+02,1.740000000000000000e+02,9.500000000000000000e+01,1.200000000000000000e+02,4.300000000000000000e+01,1.100000000000000000e+01,7.600000000000000000e+01,1.240000000000000000e+02,1.800000000000000000e+01,5.000000000000000000e+00,9.200000000000000000e+01,9.600000000000000000e+01,1.000000000000000000e+01,1.210000000000000000e+02,1.390000000000000000e+02,1.510000000000000000e+02,2.110000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.140000000000000000e+02,2.160000000000000000e+02,5.800000000000000000e+01,9.000000000000000000e+00,7.000000000000000000e+00,6.000000000000000000e+00,9.000000000000000000e+00,4.700000000000000000e+01,2.140000000000000000e+02,2.120000000000000000e+02,2.120000000000000000e+02,2.120000000000000000e+02,2.100000000000000000e+02,1.950000000000000000e+02,1.310000000000000000e+02,1.220000000000000000e+02,1.410000000000000000e+02,7.500000000000000000e+01,1.210000000000000000e+02,1.240000000000000000e+02,6.800000000000000000e+01,4.200000000000000000e+01,4.900000000000000000e+01,4.800000000000000000e+01,4.400000000000000000e+01,2.800000000000000000e+01,2.300000000000000000e+01,2.500000000000000000e+01,3.500000000000000000e+01,3.700000000000000000e+01,4.300000000000000000e+01,5.400000000000000000e+01,6.200000000000000000e+01,6.000000000000000000e+01,6.000000000000000000e+01,5.000000000000000000e+01,4.900000000000000000e+01,4.600000000000000000e+01,4.500000000000000000e+01,4.900000000000000000e+01,5.100000000000000000e+01,6.000000000000000000e+01,5.700000000000000000e+01,5.700000000000000000e+01,5.900000000000000000e+01,5.900000000000000000e+01,6.100000000000000000e+01,6.000000000000000000e+01,6.300000000000000000e+01,5.700000000000000000e+01,6.400000000000000000e+01,6.300000000000000000e+01),
(8.200000000000000000e+01,6.800000000000000000e+01,5.600000000000000000e+01,5.300000000000000000e+01,4.200000000000000000e+01,3.700000000000000000e+01,2.200000000000000000e+01,2.300000000000000000e+01,6.700000000000000000e+01,1.070000000000000000e+02,9.700000000000000000e+01,7.100000000000000000e+01,8.300000000000000000e+01,7.900000000000000000e+01,7.300000000000000000e+01,5.800000000000000000e+01,6.000000000000000000e+01,6.700000000000000000e+01,3.600000000000000000e+01,3.800000000000000000e+01,9.100000000000000000e+01,1.400000000000000000e+02,1.630000000000000000e+02,1.680000000000000000e+02,1.730000000000000000e+02,1.530000000000000000e+02,1.380000000000000000e+02,1.780000000000000000e+02,1.710000000000000000e+02,1.090000000000000000e+02,1.000000000000000000e+02,6.800000000000000000e+01,2.500000000000000000e+01,3.000000000000000000e+01,6.400000000000000000e+01,1.410000000000000000e+02,1.430000000000000000e+02,1.550000000000000000e+02,1.790000000000000000e+02,1.990000000000000000e+02,2.110000000000000000e+02,2.070000000000000000e+02,2.010000000000000000e+02,2.020000000000000000e+02,1.990000000000000000e+02,2.020000000000000000e+02,2.040000000000000000e+02,2.090000000000000000e+02,2.100000000000000000e+02,2.090000000000000000e+02,2.010000000000000000e+02,1.910000000000000000e+02,1.790000000000000000e+02,1.280000000000000000e+02,1.330000000000000000e+02,1.920000000000000000e+02,2.000000000000000000e+02,2.060000000000000000e+02,1.840000000000000000e+02,1.540000000000000000e+02,1.950000000000000000e+02,1.730000000000000000e+02,9.900000000000000000e+01,1.110000000000000000e+02,2.000000000000000000e+02,1.870000000000000000e+02,1.720000000000000000e+02,2.000000000000000000e+02,2.090000000000000000e+02,2.120000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.120000000000000000e+02,1.820000000000000000e+02,6.000000000000000000e+00,5.000000000000000000e+00,8.000000000000000000e+00,1.800000000000000000e+01,2.120000000000000000e+02,2.130000000000000000e+02,2.110000000000000000e+02,2.120000000000000000e+02,2.120000000000000000e+02,2.110000000000000000e+02,1.610000000000000000e+02,7.300000000000000000e+01,2.300000000000000000e+01,1.300000000000000000e+01,2.100000000000000000e+01,5.100000000000000000e+01,1.070000000000000000e+02,4.900000000000000000e+01,4.200000000000000000e+01,5.800000000000000000e+01,6.100000000000000000e+01,5.200000000000000000e+01,5.300000000000000000e+01,4.100000000000000000e+01,4.600000000000000000e+01,3.800000000000000000e+01,4.100000000000000000e+01,3.900000000000000000e+01,3.700000000000000000e+01,4.000000000000000000e+01,4.200000000000000000e+01,4.800000000000000000e+01,4.000000000000000000e+01,4.000000000000000000e+01,3.900000000000000000e+01,3.900000000000000000e+01,4.000000000000000000e+01,4.300000000000000000e+01,4.600000000000000000e+01,4.700000000000000000e+01,4.800000000000000000e+01,4.600000000000000000e+01,4.500000000000000000e+01,4.700000000000000000e+01,4.700000000000000000e+01,5.200000000000000000e+01,4.600000000000000000e+01,4.900000000000000000e+01,4.700000000000000000e+01),
(7.100000000000000000e+01,6.400000000000000000e+01,5.200000000000000000e+01,3.700000000000000000e+01,3.000000000000000000e+01,2.300000000000000000e+01,2.500000000000000000e+01,2.900000000000000000e+01,9.000000000000000000e+01,1.160000000000000000e+02,1.270000000000000000e+02,9.000000000000000000e+01,6.200000000000000000e+01,6.500000000000000000e+01,9.100000000000000000e+01,1.030000000000000000e+02,7.800000000000000000e+01,1.210000000000000000e+02,1.450000000000000000e+02,1.170000000000000000e+02,1.220000000000000000e+02,6.900000000000000000e+01,1.010000000000000000e+02,1.520000000000000000e+02,1.330000000000000000e+02,1.520000000000000000e+02,1.510000000000000000e+02,1.530000000000000000e+02,1.350000000000000000e+02,1.470000000000000000e+02,1.320000000000000000e+02,1.190000000000000000e+02,1.310000000000000000e+02,1.590000000000000000e+02,2.010000000000000000e+02,2.110000000000000000e+02,2.060000000000000000e+02,1.980000000000000000e+02,1.890000000000000000e+02,1.560000000000000000e+02,1.420000000000000000e+02,1.650000000000000000e+02,1.620000000000000000e+02,1.380000000000000000e+02,1.340000000000000000e+02,1.760000000000000000e+02,1.890000000000000000e+02,2.010000000000000000e+02,2.020000000000000000e+02,1.970000000000000000e+02,1.870000000000000000e+02,1.750000000000000000e+02,1.830000000000000000e+02,1.630000000000000000e+02,1.070000000000000000e+02,8.400000000000000000e+01,7.500000000000000000e+01,7.700000000000000000e+01,1.360000000000000000e+02,1.790000000000000000e+02,1.910000000000000000e+02,1.960000000000000000e+02,2.060000000000000000e+02,2.090000000000000000e+02,2.100000000000000000e+02,2.070000000000000000e+02,2.080000000000000000e+02,2.130000000000000000e+02,2.120000000000000000e+02,2.120000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.130000000000000000e+02,2.120000000000000000e+02,2.110000000000000000e+02,2.090000000000000000e+02,4.900000000000000000e+01,4.000000000000000000e+00,2.300000000000000000e+01,2.080000000000000000e+02,2.110000000000000000e+02,2.130000000000000000e+02,2.110000000000000000e+02,2.120000000000000000e+02,2.120000000000000000e+02,2.120000000000000000e+02,2.050000000000000000e+02,1.290000000000000000e+02,9.600000000000000000e+01,6.900000000000000000e+01,3.500000000000000000e+01,1.900000000000000000e+01,2.500000000000000000e+01,8.000000000000000000e+01,5.700000000000000000e+01,3.600000000000000000e+01,8.200000000000000000e+01,1.520000000000000000e+02,1.190000000000000000e+02,5.100000000000000000e+01,6.400000000000000000e+01,5.300000000000000000e+01,3.700000000000000000e+01,3.500000000000000000e+01,3.700000000000000000e+01,4.000000000000000000e+01,4.600000000000000000e+01,4.200000000000000000e+01,4.200000000000000000e+01,4.000000000000000000e+01,3.200000000000000000e+01,3.100000000000000000e+01,3.900000000000000000e+01,4.300000000000000000e+01,4.600000000000000000e+01,4.900000000000000000e+01,5.100000000000000000e+01,4.300000000000000000e+01,4.200000000000000000e+01,4.300000000000000000e+01,4.300000000000000000e+01,4.500000000000000000e+01,4.200000000000000000e+01,4.300000000000000000e+01,4.200000000000000000e+01),
(6.300000000000000000e+01,5.200000000000000000e+01,4.900000000000000000e+01,3.000000000000000000e+01,2.200000000000000000e+01,1.400000000000000000e+01,2.500000000000000000e+01,5.900000000000000000e+01,1.260000000000000000e+02,1.210000000000000000e+02,9.100000000000000000e+01,8.000000000000000000e+01,7.100000000000000000e+01,7.400000000000000000e+01,1.350000000000000000e+02,1.660000000000000000e+02,1.310000000000000000e+02,9.800000000000000000e+01,9.700000000000000000e+01,7.600000000000000000e+01,6.100000000000000000e+01,7.600000000000000000e+01,8.500000000000000000e+01,1.090000000000000000e+02,1.200000000000000000e+02,1.240000000000000000e+02,1.350000000000000000e+02,1.740000000000000000e+02,2.010000000000000000e+02,2.090000000000000000e+02,2.010000000000000000e+02,1.940000000000000000e+02,1.570000000000000000e+02,1.540000000000000000e+02,8.400000000000000000e+01,2.400000000000000000e+01,1.300000000000000000e+01,1.200000000000000000e+01,7.400000000000000000e+01,1.410000000000000000e+02,1.520000000000000000e+02,1.470000000000000000e+02,1.510000000000000000e+02,1.550000000000000000e+02,1.730000000000000000e+02,1.630000000000000000e+02,1.940000000000000000e+02,2.030000000000000000e+02,2.030000000000000000e+02,2.040000000000000000e+02,2.030000000000000000e+02,2.060000000000000000e+02,2.120000000000000000e+02,2.080000000000000000e+02,1.790000000000000000e+02,1.470000000000000000e+02,1.350000000000000000e+02,7.800000000000000000e+01,1.100000000000000000e+02,8.000000000000000000e+01,5.300000000000000000e+01,7.500000000000000000e+01,7.200000000000000000e+01,9.800000000000000000e+01,1.800000000000000000e+02,1.720000000000000000e+02,1.740000000000000000e+02,2.110000000000000000e+02,2.130000000000000000e+02,2.120000000000000000e+02,2.110000000000000000e+02,2.130000000000000000e+02,2.120000000000000000e+02,2.100000000000000000e+02,2.110000000000000000e+02,2.100000000000000000e+02,1.960000000000000000e+02,2.010000000000000000e+02,1.970000000000000000e+02,1.290000000000000000e+02,8.000000000000000000e+00,1.810000000000000000e+02,2.120000000000000000e+02,2.110000000000000000e+02,2.110000000000000000e+02,2.130000000000000000e+02,2.110000000000000000e+02,2.110000000000000000e+02,2.090000000000000000e+02,2.080000000000000000e+02,2.060000000000000000e+02,1.820000000000000000e+02,1.820000000000000000e+02,1.370000000000000000e+02,1.060000000000000000e+02,9.000000000000000000e+01,2.500000000000000000e+01,1.300000000000000000e+01,4.000000000000000000e+01,8.700000000000000000e+01,8.800000000000000000e+01,6.300000000000000000e+01,1.040000000000000000e+02,1.660000000000000000e+02,1.510000000000000000e+02,9.600000000000000000e+01,5.800000000000000000e+01,3.700000000000000000e+01,4.500000000000000000e+01,4.800000000000000000e+01,3.700000000000000000e+01,4.000000000000000000e+01,4.400000000000000000e+01,3.900000000000000000e+01,4.200000000000000000e+01,3.700000000000000000e+01,3.200000000000000000e+01,3.900000000000000000e+01,4.600000000000000000e+01,5.100000000000000000e+01,4.400000000000000000e+01,4.500000000000000000e+01,4.400000000000000000e+01,4.600000000000000000e+01,4.600000000000000000e+01,4.000000000000000000e+01,4.400000000000000000e+01,4.000000000000000000e+01),
(5.400000000000000000e+01,4.000000000000000000e+01,3.400000000000000000e+01,2.400000000000000000e+01,1.700000000000000000e+01,1.500000000000000000e+01,3.700000000000000000e+01,1.080000000000000000e+02,1.480000000000000000e+02,1.400000000000000000e+02,1.070000000000000000e+02,6.000000000000000000e+01,1.040000000000000000e+02,1.300000000000000000e+02,1.060000000000000000e+02,1.270000000000000000e+02,1.090000000000000000e+02,1.010000000000000000e+02,6.000000000000000000e+01,1.140000000000000000e+02,1.110000000000000000e+02,4.700000000000000000e+01,3.300000000000000000e+01,6.500000000000000000e+01,1.530000000000000000e+02,2.010000000000000000e+02,2.110000000000000000e+02,2.020000000000000000e+02,1.760000000000000000e+02,1.760000000000000000e+02,1.840000000000000000e+02,1.740000000000000000e+02,1.440000000000000000e+02,1.190000000000000000e+02,8.700000000000000000e+01,7.000000000000000000e+01,7.500000000000000000e+01,7.400000000000000000e+01,7.900000000000000000e+01,9.200000000000000000e+01,1.480000000000000000e+02,1.400000000000000000e+02,1.270000000000000000e+02,1.450000000000000000e+02,1.580000000000000000e+02,1.900000000000000000e+02,2.090000000000000000e+02,2.120000000000000000e+02,2.120000000000000000e+02,2.090000000000000000e+02,2.020000000000000000e+02,1.890000000000000000e+02,1.910000000000000000e+02,1.240000000000000000e+02,4.000000000000000000e+01,9.000000000000000000e+01,1.950000000000000000e+02,1.920000000000000000e+02,1.670000000000000000e+02,1.500000000000000000e+02,1.570000000000000000e+02,1.980000000000000000e+02,1.590000000000000000e+02,1.350000000000000000e+02,2.090000000000000000e+02,2.080000000000000000e+02,2.010000000000000000e+02,2.070000000000000000e+02,2.120000000000000000e+02,2.040000000000000000e+02,2.080000000000000000e+02,2.130000000000000000e+02,2.110000000000000000e+02,1.990000000000000000e+02,2.080000000000000000e+02,2.070000000000000000e+02,1.990000000000000000e+02,2.060000000000000000e+02,1.740000000000000000e+02,1.080000000000000000e+02,5.500000000000000000e+01,1.900000000000000000e+02,2.020000000000000000e+02,2.120000000000000000e+02,2.060000000000000000e+02,2.100000000000000000e+02,2.090000000000000000e+02,2.090000000000000000e+02,2.090000000000000000e+02,1.980000000000000000e+02,1.970000000000000000e+02,1.730000000000000000e+02,1.660000000000000000e+02,1.260000000000000000e+02,8.000000000000000000e+01,5.200000000000000000e+01,2.900000000000000000e+01,4.200000000000000000e+01,6.900000000000000000e+01,1.400000000000000000e+02,1.470000000000000000e+02,7.800000000000000000e+01,9.100000000000000000e+01,6.700000000000000000e+01,3.800000000000000000e+01,5.100000000000000000e+01,8.500000000000000000e+01,1.210000000000000000e+02,9.700000000000000000e+01,5.500000000000000000e+01,4.500000000000000000e+01,4.100000000000000000e+01,3.900000000000000000e+01,3.500000000000000000e+01,3.900000000000000000e+01,4.300000000000000000e+01,4.100000000000000000e+01,3.600000000000000000e+01,4.600000000000000000e+01,5.000000000000000000e+01,4.500000000000000000e+01,5.100000000000000000e+01,4.400000000000000000e+01,4.200000000000000000e+01,4.300000000000000000e+01,4.300000000000000000e+01,4.400000000000000000e+01,4.100000000000000000e+01),
(4.800000000000000000e+01,3.200000000000000000e+01,2.200000000000000000e+01,2.000000000000000000e+01,1.700000000000000000e+01,3.600000000000000000e+01,4.700000000000000000e+01,1.050000000000000000e+02,1.430000000000000000e+02,1.370000000000000000e+02,1.180000000000000000e+02,9.800000000000000000e+01,5.100000000000000000e+01,6.900000000000000000e+01,1.250000000000000000e+02,1.230000000000000000e+02,1.140000000000000000e+02,1.110000000000000000e+02,4.800000000000000000e+01,8.300000000000000000e+01,9.300000000000000000e+01,8.600000000000000000e+01,1.400000000000000000e+02,1.720000000000000000e+02,1.140000000000000000e+02,1.010000000000000000e+02,1.550000000000000000e+02,1.690000000000000000e+02,1.750000000000000000e+02,1.750000000000000000e+02,1.610000000000000000e+02,1.580000000000000000e+02,1.330000000000000000e+02,1.090000000000000000e+02,9.700000000000000000e+01,7.100000000000000000e+01,4.000000000000000000e+01,4.100000000000000000e+01,2.200000000000000000e+01,1.600000000000000000e+01,3.800000000000000000e+01,1.360000000000000000e+02,2.020000000000000000e+02,2.120000000000000000e+02,2.080000000000000000e+02,2.000000000000000000e+02,2.040000000000000000e+02,2.000000000000000000e+02,1.960000000000000000e+02,1.980000000000000000e+02,1.980000000000000000e+02,2.010000000000000000e+02,1.940000000000000000e+02,2.010000000000000000e+02,1.800000000000000000e+02,1.430000000000000000e+02,1.340000000000000000e+02,8.300000000000000000e+01,1.030000000000000000e+02,1.060000000000000000e+02,1.650000000000000000e+02,1.910000000000000000e+02,1.990000000000000000e+02,2.070000000000000000e+02,2.120000000000000000e+02,2.120000000000000000e+02,2.120000000000000000e+02,2.120000000000000000e+02,2.140000000000000000e+02,2.130000000000000000e+02,2.110000000000000000e+02,2.130000000000000000e+02,2.120000000000000000e+02,2.120000000000000000e+02,2.140000000000000000e+02,1.830000000000000000e+02,1.990000000000000000e+02,1.270000000000000000e+02,9.200000000000000000e+01,4.400000000000000000e+01,1.110000000000000000e+02,1.800000000000000000e+02,2.080000000000000000e+02,2.130000000000000000e+02,2.080000000000000000e+02,2.100000000000000000e+02,1.950000000000000000e+02,1.970000000000000000e+02,1.900000000000000000e+02,1.580000000000000000e+02,1.490000000000000000e+02,9.300000000000000000e+01,3.100000000000000000e+01,2.600000000000000000e+01,3.800000000000000000e+01,5.800000000000000000e+01,2.600000000000000000e+01,1.900000000000000000e+01,2.800000000000000000e+01,3.000000000000000000e+01,5.300000000000000000e+01,1.280000000000000000e+02,1.780000000000000000e+02,1.010000000000000000e+02,4.000000000000000000e+01,3.300000000000000000e+01,3.200000000000000000e+01,3.300000000000000000e+01,3.700000000000000000e+01,6.300000000000000000e+01,9.500000000000000000e+01,9.900000000000000000e+01,5.800000000000000000e+01,3.000000000000000000e+01,3.200000000000000000e+01,3.300000000000000000e+01,3.300000000000000000e+01,3.600000000000000000e+01,3.700000000000000000e+01,3.400000000000000000e+01,4.000000000000000000e+01,4.000000000000000000e+01,3.900000000000000000e+01,3.900000000000000000e+01,3.400000000000000000e+01,3.400000000000000000e+01,3.500000000000000000e+01,3.300000000000000000e+01),
(3.900000000000000000e+01,3.800000000000000000e+01,2.200000000000000000e+01,3.200000000000000000e+01,3.500000000000000000e+01,3.000000000000000000e+01,8.000000000000000000e+01,1.130000000000000000e+02,1.300000000000000000e+02,1.170000000000000000e+02,7.900000000000000000e+01,9.800000000000000000e+01,9.100000000000000000e+01,8.000000000000000000e+01,8.700000000000000000e+01,8.800000000000000000e+01,1.080000000000000000e+02,8.500000000000000000e+01,5.000000000000000000e+01,6.000000000000000000e+01,1.530000000000000000e+02,1.700000000000000000e+02,9.600000000000000000e+01,4.800000000000000000e+01,7.400000000000000000e+01,8.500000000000000000e+01,1.060000000000000000e+02,1.740000000000000000e+02,1.360000000000000000e+02,1.220000000000000000e+02,1.370000000000000000e+02,1.230000000000000000e+02,1.440000000000000000e+02,1.530000000000000000e+02,1.110000000000000000e+02,5.500000000000000000e+01,3.600000000000000000e+01,2.400000000000000000e+01,1.210000000000000000e+02,2.060000000000000000e+02,1.520000000000000000e+02,1.240000000000000000e+02,6.300000000000000000e+01,1.030000000000000000e+02,1.520000000000000000e+02,1.610000000000000000e+02,1.830000000000000000e+02,1.890000000000000000e+02,1.860000000000000000e+02,2.080000000000000000e+02,2.090000000000000000e+02,2.070000000000000000e+02,2.080000000000000000e+02,1.990000000000000000e+02,1.850000000000000000e+02,1.010000000000000000e+02,1.060000000000000000e+02,1.000000000000000000e+02,1.040000000000000000e+02,1.280000000000000000e+02,1.150000000000000000e+02,1.050000000000000000e+02,1.320000000000000000e+02,1.800000000000000000e+02,1.680000000000000000e+02,2.090000000000000000e+02,2.080000000000000000e+02,2.080000000000000000e+02,2.070000000000000000e+02,2.110000000000000000e+02,2.130000000000000000e+02,2.110000000000000000e+02,2.110000000000000000e+02,2.110000000000000000e+02,2.150000000000000000e+02,1.790000000000000000e+02,1.700000000000000000e+02,1.450000000000000000e+02,6.700000000000000000e+01,2.300000000000000000e+01,7.500000000000000000e+01,1.320000000000000000e+02,2.080000000000000000e+02,1.870000000000000000e+02,2.100000000000000000e+02,2.080000000000000000e+02,2.040000000000000000e+02,2.120000000000000000e+02,1.940000000000000000e+02,2.010000000000000000e+02,1.990000000000000000e+02,1.520000000000000000e+02,1.480000000000000000e+02,1.500000000000000000e+02,1.430000000000000000e+02,1.460000000000000000e+02,1.490000000000000000e+02,2.800000000000000000e+01,2.400000000000000000e+01,3.700000000000000000e+01,5.500000000000000000e+01,9.100000000000000000e+01,9.400000000000000000e+01,1.070000000000000000e+02,1.120000000000000000e+02,2.500000000000000000e+01,1.800000000000000000e+01,1.700000000000000000e+01,2.000000000000000000e+01,1.900000000000000000e+01,1.800000000000000000e+01,1.900000000000000000e+01,4.900000000000000000e+01,6.700000000000000000e+01,4.200000000000000000e+01,2.100000000000000000e+01,2.000000000000000000e+01,2.000000000000000000e+01,1.900000000000000000e+01,1.900000000000000000e+01,1.800000000000000000e+01,1.800000000000000000e+01,2.100000000000000000e+01,2.100000000000000000e+01,2.100000000000000000e+01,2.100000000000000000e+01,2.200000000000000000e+01,1.900000000000000000e+01),
(4.800000000000000000e+01,4.300000000000000000e+01,4.400000000000000000e+01,3.500000000000000000e+01,2.800000000000000000e+01,4.400000000000000000e+01,1.110000000000000000e+02,1.420000000000000000e+02,1.460000000000000000e+02,1.110000000000000000e+02,8.000000000000000000e+01,8.700000000000000000e+01,8.500000000000000000e+01,6.800000000000000000e+01,1.050000000000000000e+02,7.900000000000000000e+01,8.900000000000000000e+01,7.500000000000000000e+01,1.400000000000000000e+02,8.200000000000000000e+01,1.270000000000000000e+02,1.240000000000000000e+02,1.380000000000000000e+02,1.020000000000000000e+02,7.500000000000000000e+01,8.900000000000000000e+01,1.490000000000000000e+02,1.290000000000000000e+02,1.640000000000000000e+02,1.780000000000000000e+02,1.640000000000000000e+02,1.610000000000000000e+02,1.370000000000000000e+02,1.640000000000000000e+02,1.500000000000000000e+02,1.910000000000000000e+02,1.850000000000000000e+02,1.090000000000000000e+02,1.000000000000000000e+01,2.600000000000000000e+01,1.900000000000000000e+01,1.500000000000000000e+01,1.200000000000000000e+01,4.000000000000000000e+01,1.200000000000000000e+02,1.590000000000000000e+02,1.630000000000000000e+02,1.900000000000000000e+02,2.110000000000000000e+02,2.090000000000000000e+02,2.070000000000000000e+02,2.070000000000000000e+02,2.070000000000000000e+02,2.010000000000000000e+02,1.870000000000000000e+02,1.680000000000000000e+02,1.360000000000000000e+02,1.220000000000000000e+02,5.000000000000000000e+01,9.000000000000000000e+01,7.900000000000000000e+01,1.340000000000000000e+02,1.830000000000000000e+02,1.690000000000000000e+02,1.960000000000000000e+02,1.980000000000000000e+02,2.030000000000000000e+02,2.050000000000000000e+02,2.100000000000000000e+02,2.120000000000000000e+02,2.110000000000000000e+02,2.070000000000000000e+02,2.040000000000000000e+02,2.090000000000000000e+02,1.730000000000000000e+02,1.770000000000000000e+02,1.000000000000000000e+02,1.210000000000000000e+02,5.800000000000000000e+01,5.700000000000000000e+01,7.800000000000000000e+01,1.090000000000000000e+02,1.870000000000000000e+02,2.040000000000000000e+02,1.990000000000000000e+02,1.990000000000000000e+02,2.040000000000000000e+02,2.100000000000000000e+02,2.040000000000000000e+02,1.950000000000000000e+02,1.890000000000000000e+02,1.650000000000000000e+02,9.400000000000000000e+01,4.900000000000000000e+01,1.320000000000000000e+02,1.390000000000000000e+02,9.600000000000000000e+01,1.340000000000000000e+02,1.580000000000000000e+02,1.040000000000000000e+02,1.040000000000000000e+02,1.220000000000000000e+02,8.700000000000000000e+01,2.300000000000000000e+01,1.400000000000000000e+01,5.100000000000000000e+01,8.400000000000000000e+01,1.100000000000000000e+01,7.000000000000000000e+00,6.000000000000000000e+00,6.000000000000000000e+00,8.000000000000000000e+00,7.000000000000000000e+00,9.000000000000000000e+00,1.700000000000000000e+01,4.000000000000000000e+01,1.400000000000000000e+01,7.000000000000000000e+00,9.000000000000000000e+00,9.000000000000000000e+00,7.000000000000000000e+00,7.000000000000000000e+00,8.000000000000000000e+00,9.000000000000000000e+00,1.000000000000000000e+01,1.000000000000000000e+01,8.000000000000000000e+00,1.000000000000000000e+01),
(4.900000000000000000e+01,6.000000000000000000e+01,2.600000000000000000e+01,3.800000000000000000e+01,5.100000000000000000e+01,6.900000000000000000e+01,1.470000000000000000e+02,1.610000000000000000e+02,1.390000000000000000e+02,1.240000000000000000e+02,9.100000000000000000e+01,6.800000000000000000e+01,1.160000000000000000e+02,1.200000000000000000e+02,1.250000000000000000e+02,1.240000000000000000e+02,1.450000000000000000e+02,8.800000000000000000e+01,3.800000000000000000e+01,4.000000000000000000e+01,4.900000000000000000e+01,1.020000000000000000e+02,9.200000000000000000e+01,1.090000000000000000e+02,1.620000000000000000e+02,1.290000000000000000e+02,9.700000000000000000e+01,1.450000000000000000e+02,1.790000000000000000e+02,1.600000000000000000e+02,1.360000000000000000e+02,1.630000000000000000e+02,2.030000000000000000e+02,1.930000000000000000e+02,1.660000000000000000e+02,1.510000000000000000e+02,7.600000000000000000e+01,3.400000000000000000e+01,1.900000000000000000e+01,1.200000000000000000e+01,1.000000000000000000e+01,2.300000000000000000e+01,3.000000000000000000e+01,2.900000000000000000e+01,6.000000000000000000e+01,1.770000000000000000e+02,1.810000000000000000e+02,1.920000000000000000e+02,1.670000000000000000e+02,1.830000000000000000e+02,2.030000000000000000e+02,2.050000000000000000e+02,2.060000000000000000e+02,2.030000000000000000e+02,2.040000000000000000e+02,1.980000000000000000e+02,1.960000000000000000e+02,1.320000000000000000e+02,1.290000000000000000e+02,9.000000000000000000e+01,1.170000000000000000e+02,6.100000000000000000e+01,1.510000000000000000e+02,1.780000000000000000e+02,1.730000000000000000e+02,1.880000000000000000e+02,2.010000000000000000e+02,2.070000000000000000e+02,2.080000000000000000e+02,1.950000000000000000e+02,2.050000000000000000e+02,1.980000000000000000e+02,1.810000000000000000e+02,1.380000000000000000e+02,1.260000000000000000e+02,1.500000000000000000e+02,1.370000000000000000e+02,1.230000000000000000e+02,1.460000000000000000e+02,1.520000000000000000e+02,1.400000000000000000e+02,1.240000000000000000e+02,1.320000000000000000e+02,1.790000000000000000e+02,1.830000000000000000e+02,1.910000000000000000e+02,1.970000000000000000e+02,1.880000000000000000e+02,1.410000000000000000e+02,1.070000000000000000e+02,9.800000000000000000e+01,7.400000000000000000e+01,5.600000000000000000e+01,2.500000000000000000e+01,1.500000000000000000e+01,5.800000000000000000e+01,9.400000000000000000e+01,1.750000000000000000e+02,1.330000000000000000e+02,1.760000000000000000e+02,1.660000000000000000e+02,9.500000000000000000e+01,7.500000000000000000e+01,3.200000000000000000e+01,2.500000000000000000e+01,1.700000000000000000e+01,1.500000000000000000e+01,5.400000000000000000e+01,6.700000000000000000e+01,1.200000000000000000e+01,1.200000000000000000e+01,1.400000000000000000e+01,1.300000000000000000e+01,1.500000000000000000e+01,1.500000000000000000e+01,1.200000000000000000e+01,2.900000000000000000e+01,3.000000000000000000e+01,1.300000000000000000e+01,1.300000000000000000e+01,1.300000000000000000e+01,1.600000000000000000e+01,1.600000000000000000e+01,1.500000000000000000e+01,1.700000000000000000e+01,1.700000000000000000e+01,1.600000000000000000e+01,1.800000000000000000e+01),
(6.200000000000000000e+01,4.900000000000000000e+01,3.300000000000000000e+01,4.400000000000000000e+01,7.600000000000000000e+01,1.070000000000000000e+02,1.250000000000000000e+02,1.690000000000000000e+02,1.550000000000000000e+02,1.300000000000000000e+02,1.210000000000000000e+02,7.900000000000000000e+01,7.400000000000000000e+01,9.900000000000000000e+01,1.090000000000000000e+02,1.510000000000000000e+02,8.700000000000000000e+01,6.200000000000000000e+01,4.400000000000000000e+01,2.100000000000000000e+01,4.300000000000000000e+01,8.100000000000000000e+01,1.280000000000000000e+02,1.570000000000000000e+02,8.300000000000000000e+01,7.800000000000000000e+01,9.700000000000000000e+01,1.210000000000000000e+02,1.610000000000000000e+02,1.620000000000000000e+02,1.940000000000000000e+02,1.480000000000000000e+02,1.580000000000000000e+02,1.710000000000000000e+02,1.800000000000000000e+02,1.360000000000000000e+02,1.040000000000000000e+02,9.400000000000000000e+01,7.100000000000000000e+01,4.000000000000000000e+01,3.000000000000000000e+01,1.900000000000000000e+01,2.100000000000000000e+01,1.210000000000000000e+02,7.700000000000000000e+01,1.610000000000000000e+02,1.030000000000000000e+02,1.030000000000000000e+02,1.240000000000000000e+02,1.520000000000000000e+02,1.770000000000000000e+02,2.050000000000000000e+02,2.000000000000000000e+02,2.050000000000000000e+02,2.070000000000000000e+02,1.990000000000000000e+02,1.850000000000000000e+02,1.960000000000000000e+02,1.850000000000000000e+02,1.740000000000000000e+02,8.600000000000000000e+01,1.200000000000000000e+02,1.590000000000000000e+02,1.330000000000000000e+02,1.800000000000000000e+02,1.920000000000000000e+02,1.970000000000000000e+02,1.850000000000000000e+02,1.640000000000000000e+02,1.520000000000000000e+02,1.610000000000000000e+02,1.600000000000000000e+02,1.710000000000000000e+02,1.660000000000000000e+02,1.760000000000000000e+02,1.640000000000000000e+02,1.890000000000000000e+02,1.880000000000000000e+02,1.940000000000000000e+02,2.040000000000000000e+02,1.880000000000000000e+02,1.600000000000000000e+02,1.380000000000000000e+02,1.240000000000000000e+02,1.380000000000000000e+02,1.840000000000000000e+02,1.900000000000000000e+02,1.890000000000000000e+02,1.840000000000000000e+02,1.570000000000000000e+02,6.200000000000000000e+01,2.900000000000000000e+01,3.900000000000000000e+01,7.500000000000000000e+01,3.700000000000000000e+01,3.500000000000000000e+01,9.700000000000000000e+01,1.370000000000000000e+02,1.660000000000000000e+02,1.650000000000000000e+02,1.150000000000000000e+02,1.760000000000000000e+02,9.900000000000000000e+01,6.000000000000000000e+01,4.200000000000000000e+01,4.700000000000000000e+01,4.000000000000000000e+01,3.800000000000000000e+01,5.300000000000000000e+01,1.070000000000000000e+02,4.600000000000000000e+01,4.000000000000000000e+01,3.900000000000000000e+01,3.800000000000000000e+01,4.000000000000000000e+01,4.300000000000000000e+01,4.600000000000000000e+01,5.800000000000000000e+01,4.800000000000000000e+01,4.500000000000000000e+01,4.600000000000000000e+01,4.400000000000000000e+01,4.600000000000000000e+01,4.500000000000000000e+01,4.200000000000000000e+01,4.200000000000000000e+01,4.800000000000000000e+01,5.000000000000000000e+01),
(6.200000000000000000e+01,5.500000000000000000e+01,4.700000000000000000e+01,8.000000000000000000e+01,1.250000000000000000e+02,1.200000000000000000e+02,1.180000000000000000e+02,1.280000000000000000e+02,1.350000000000000000e+02,1.120000000000000000e+02,1.020000000000000000e+02,7.100000000000000000e+01,9.200000000000000000e+01,1.410000000000000000e+02,1.290000000000000000e+02,9.800000000000000000e+01,7.300000000000000000e+01,7.600000000000000000e+01,4.200000000000000000e+01,2.100000000000000000e+01,2.000000000000000000e+01,7.900000000000000000e+01,1.430000000000000000e+02,1.170000000000000000e+02,9.900000000000000000e+01,8.800000000000000000e+01,6.600000000000000000e+01,1.040000000000000000e+02,1.660000000000000000e+02,1.520000000000000000e+02,1.710000000000000000e+02,1.750000000000000000e+02,1.870000000000000000e+02,1.790000000000000000e+02,1.670000000000000000e+02,1.200000000000000000e+02,1.010000000000000000e+02,1.000000000000000000e+02,1.040000000000000000e+02,9.800000000000000000e+01,6.900000000000000000e+01,1.130000000000000000e+02,5.700000000000000000e+01,7.800000000000000000e+01,4.000000000000000000e+01,2.100000000000000000e+01,5.900000000000000000e+01,1.040000000000000000e+02,8.600000000000000000e+01,1.330000000000000000e+02,1.560000000000000000e+02,1.590000000000000000e+02,1.920000000000000000e+02,2.040000000000000000e+02,1.930000000000000000e+02,2.020000000000000000e+02,2.030000000000000000e+02,2.090000000000000000e+02,2.020000000000000000e+02,1.580000000000000000e+02,1.720000000000000000e+02,1.980000000000000000e+02,1.710000000000000000e+02,1.590000000000000000e+02,1.560000000000000000e+02,1.870000000000000000e+02,1.730000000000000000e+02,1.420000000000000000e+02,1.660000000000000000e+02,1.860000000000000000e+02,1.990000000000000000e+02,1.960000000000000000e+02,2.040000000000000000e+02,2.010000000000000000e+02,2.100000000000000000e+02,2.070000000000000000e+02,2.080000000000000000e+02,2.030000000000000000e+02,2.090000000000000000e+02,2.090000000000000000e+02,2.060000000000000000e+02,1.830000000000000000e+02,1.850000000000000000e+02,1.600000000000000000e+02,9.100000000000000000e+01,1.480000000000000000e+02,1.620000000000000000e+02,1.410000000000000000e+02,8.400000000000000000e+01,1.000000000000000000e+02,4.700000000000000000e+01,3.100000000000000000e+01,9.000000000000000000e+00,1.200000000000000000e+01,1.110000000000000000e+02,1.030000000000000000e+02,1.000000000000000000e+02,1.480000000000000000e+02,1.620000000000000000e+02,1.710000000000000000e+02,1.600000000000000000e+02,1.440000000000000000e+02,1.410000000000000000e+02,9.700000000000000000e+01,7.800000000000000000e+01,9.000000000000000000e+01,8.500000000000000000e+01,7.300000000000000000e+01,6.700000000000000000e+01,6.600000000000000000e+01,1.090000000000000000e+02,1.010000000000000000e+02,6.300000000000000000e+01,6.900000000000000000e+01,6.500000000000000000e+01,7.100000000000000000e+01,6.700000000000000000e+01,7.200000000000000000e+01,7.900000000000000000e+01,7.600000000000000000e+01,7.000000000000000000e+01,7.600000000000000000e+01,7.700000000000000000e+01,7.600000000000000000e+01,7.500000000000000000e+01,7.600000000000000000e+01,7.800000000000000000e+01,7.300000000000000000e+01),
(5.300000000000000000e+01,5.800000000000000000e+01,5.400000000000000000e+01,8.000000000000000000e+01,1.110000000000000000e+02,1.190000000000000000e+02,1.090000000000000000e+02,1.140000000000000000e+02,1.040000000000000000e+02,1.020000000000000000e+02,9.400000000000000000e+01,8.600000000000000000e+01,1.170000000000000000e+02,9.800000000000000000e+01,1.630000000000000000e+02,1.380000000000000000e+02,8.500000000000000000e+01,5.800000000000000000e+01,3.700000000000000000e+01,2.300000000000000000e+01,2.600000000000000000e+01,9.400000000000000000e+01,8.900000000000000000e+01,1.110000000000000000e+02,1.080000000000000000e+02,1.120000000000000000e+02,1.850000000000000000e+02,1.190000000000000000e+02,9.100000000000000000e+01,1.310000000000000000e+02,1.430000000000000000e+02,1.840000000000000000e+02,1.780000000000000000e+02,1.510000000000000000e+02,1.100000000000000000e+02,1.240000000000000000e+02,1.260000000000000000e+02,1.830000000000000000e+02,1.510000000000000000e+02,1.710000000000000000e+02,1.890000000000000000e+02,1.520000000000000000e+02,1.550000000000000000e+02,5.500000000000000000e+01,3.600000000000000000e+01,1.500000000000000000e+01,2.000000000000000000e+01,6.400000000000000000e+01,7.400000000000000000e+01,5.900000000000000000e+01,1.640000000000000000e+02,1.660000000000000000e+02,1.840000000000000000e+02,2.030000000000000000e+02,1.680000000000000000e+02,2.010000000000000000e+02,2.030000000000000000e+02,2.070000000000000000e+02,2.000000000000000000e+02,1.890000000000000000e+02,2.060000000000000000e+02,1.950000000000000000e+02,1.930000000000000000e+02,1.810000000000000000e+02,1.710000000000000000e+02,2.080000000000000000e+02,2.050000000000000000e+02,2.050000000000000000e+02,2.070000000000000000e+02,2.080000000000000000e+02,2.070000000000000000e+02,2.100000000000000000e+02,2.090000000000000000e+02,2.090000000000000000e+02,2.100000000000000000e+02,2.100000000000000000e+02,2.070000000000000000e+02,2.100000000000000000e+02,2.090000000000000000e+02,2.090000000000000000e+02,2.100000000000000000e+02,2.090000000000000000e+02,2.080000000000000000e+02,1.980000000000000000e+02,1.530000000000000000e+02,1.140000000000000000e+02,1.050000000000000000e+02,1.050000000000000000e+02,5.200000000000000000e+01,3.300000000000000000e+01,2.500000000000000000e+01,3.000000000000000000e+01,6.000000000000000000e+01,3.100000000000000000e+01,6.000000000000000000e+01,1.310000000000000000e+02,1.430000000000000000e+02,1.570000000000000000e+02,1.410000000000000000e+02,1.520000000000000000e+02,1.380000000000000000e+02,8.400000000000000000e+01,1.120000000000000000e+02,1.260000000000000000e+02,1.440000000000000000e+02,1.200000000000000000e+02,1.140000000000000000e+02,1.380000000000000000e+02,1.420000000000000000e+02,1.340000000000000000e+02,1.300000000000000000e+02,1.400000000000000000e+02,1.570000000000000000e+02,1.290000000000000000e+02,1.320000000000000000e+02,1.340000000000000000e+02,1.330000000000000000e+02,1.340000000000000000e+02,1.370000000000000000e+02,1.400000000000000000e+02,1.330000000000000000e+02,1.370000000000000000e+02,1.380000000000000000e+02,1.410000000000000000e+02,1.330000000000000000e+02,1.300000000000000000e+02,1.370000000000000000e+02,1.370000000000000000e+02),
(5.900000000000000000e+01,4.600000000000000000e+01,4.900000000000000000e+01,9.700000000000000000e+01,1.020000000000000000e+02,1.100000000000000000e+02,1.160000000000000000e+02,1.100000000000000000e+02,1.310000000000000000e+02,1.390000000000000000e+02,1.380000000000000000e+02,1.190000000000000000e+02,7.000000000000000000e+01,1.180000000000000000e+02,1.100000000000000000e+02,1.330000000000000000e+02,9.400000000000000000e+01,6.900000000000000000e+01,5.400000000000000000e+01,5.600000000000000000e+01,8.700000000000000000e+01,3.800000000000000000e+01,4.200000000000000000e+01,1.020000000000000000e+02,1.310000000000000000e+02,1.770000000000000000e+02,1.330000000000000000e+02,1.130000000000000000e+02,9.200000000000000000e+01,1.090000000000000000e+02,1.450000000000000000e+02,1.730000000000000000e+02,1.940000000000000000e+02,2.020000000000000000e+02,2.020000000000000000e+02,1.970000000000000000e+02,1.730000000000000000e+02,1.690000000000000000e+02,1.990000000000000000e+02,1.750000000000000000e+02,1.800000000000000000e+02,1.780000000000000000e+02,1.280000000000000000e+02,8.300000000000000000e+01,8.200000000000000000e+01,3.700000000000000000e+01,3.200000000000000000e+01,3.100000000000000000e+01,1.380000000000000000e+02,2.010000000000000000e+02,1.580000000000000000e+02,1.690000000000000000e+02,1.630000000000000000e+02,1.910000000000000000e+02,1.480000000000000000e+02,2.020000000000000000e+02,1.730000000000000000e+02,2.070000000000000000e+02,1.980000000000000000e+02,2.030000000000000000e+02,1.880000000000000000e+02,1.950000000000000000e+02,1.970000000000000000e+02,1.970000000000000000e+02,2.070000000000000000e+02,2.100000000000000000e+02,2.090000000000000000e+02,2.100000000000000000e+02,2.100000000000000000e+02,2.120000000000000000e+02,2.120000000000000000e+02,2.120000000000000000e+02,2.120000000000000000e+02,2.120000000000000000e+02,2.100000000000000000e+02,2.100000000000000000e+02,2.090000000000000000e+02,2.060000000000000000e+02,2.110000000000000000e+02,2.110000000000000000e+02,2.110000000000000000e+02,2.100000000000000000e+02,2.130000000000000000e+02,2.070000000000000000e+02,1.890000000000000000e+02,1.800000000000000000e+02,1.090000000000000000e+02,6.600000000000000000e+01,4.500000000000000000e+01,4.400000000000000000e+01,9.700000000000000000e+01,4.200000000000000000e+01,4.500000000000000000e+01,9.700000000000000000e+01,1.040000000000000000e+02,1.200000000000000000e+02,1.590000000000000000e+02,1.440000000000000000e+02,1.460000000000000000e+02,1.160000000000000000e+02,9.500000000000000000e+01,7.600000000000000000e+01,7.800000000000000000e+01,1.460000000000000000e+02,1.680000000000000000e+02,1.810000000000000000e+02,1.670000000000000000e+02,1.690000000000000000e+02,1.800000000000000000e+02,1.810000000000000000e+02,1.810000000000000000e+02,1.800000000000000000e+02,1.820000000000000000e+02,1.890000000000000000e+02,1.830000000000000000e+02,1.780000000000000000e+02,1.810000000000000000e+02,1.820000000000000000e+02,1.820000000000000000e+02,1.860000000000000000e+02,1.780000000000000000e+02,1.790000000000000000e+02,1.820000000000000000e+02,1.850000000000000000e+02,1.820000000000000000e+02,1.820000000000000000e+02,1.800000000000000000e+02,1.830000000000000000e+02),
(5.800000000000000000e+01,4.100000000000000000e+01,7.000000000000000000e+01,1.130000000000000000e+02,1.180000000000000000e+02,1.100000000000000000e+02,7.900000000000000000e+01,7.700000000000000000e+01,1.000000000000000000e+02,1.160000000000000000e+02,1.010000000000000000e+02,1.150000000000000000e+02,8.500000000000000000e+01,9.900000000000000000e+01,1.590000000000000000e+02,1.460000000000000000e+02,5.900000000000000000e+01,3.100000000000000000e+01,3.300000000000000000e+01,5.800000000000000000e+01,3.500000000000000000e+01,4.800000000000000000e+01,8.900000000000000000e+01,1.230000000000000000e+02,1.280000000000000000e+02,1.180000000000000000e+02,1.350000000000000000e+02,1.360000000000000000e+02,7.900000000000000000e+01,1.440000000000000000e+02,1.660000000000000000e+02,1.790000000000000000e+02,1.720000000000000000e+02,1.670000000000000000e+02,1.830000000000000000e+02,1.890000000000000000e+02,1.880000000000000000e+02,1.990000000000000000e+02,1.840000000000000000e+02,1.720000000000000000e+02,1.750000000000000000e+02,1.610000000000000000e+02,1.670000000000000000e+02,1.560000000000000000e+02,1.230000000000000000e+02,9.700000000000000000e+01,6.200000000000000000e+01,7.000000000000000000e+01,4.800000000000000000e+01,5.700000000000000000e+01,9.700000000000000000e+01,1.460000000000000000e+02,1.600000000000000000e+02,1.690000000000000000e+02,1.790000000000000000e+02,1.600000000000000000e+02,1.850000000000000000e+02,2.020000000000000000e+02,1.930000000000000000e+02,2.020000000000000000e+02,1.760000000000000000e+02,2.010000000000000000e+02,1.920000000000000000e+02,2.020000000000000000e+02,2.080000000000000000e+02,2.090000000000000000e+02,2.090000000000000000e+02,2.110000000000000000e+02,2.110000000000000000e+02,2.120000000000000000e+02,2.100000000000000000e+02,2.080000000000000000e+02,2.110000000000000000e+02,2.110000000000000000e+02,2.100000000000000000e+02,2.080000000000000000e+02,2.100000000000000000e+02,2.080000000000000000e+02,2.090000000000000000e+02,2.100000000000000000e+02,2.130000000000000000e+02,2.120000000000000000e+02,2.090000000000000000e+02,2.080000000000000000e+02,1.860000000000000000e+02,1.330000000000000000e+02,1.090000000000000000e+02,5.500000000000000000e+01,2.700000000000000000e+01,1.000000000000000000e+01,3.000000000000000000e+01,3.200000000000000000e+01,9.700000000000000000e+01,1.270000000000000000e+02,1.320000000000000000e+02,1.450000000000000000e+02,1.530000000000000000e+02,1.710000000000000000e+02,1.030000000000000000e+02,6.400000000000000000e+01,5.800000000000000000e+01,4.100000000000000000e+01,6.900000000000000000e+01,1.460000000000000000e+02,1.850000000000000000e+02,1.890000000000000000e+02,1.920000000000000000e+02,1.930000000000000000e+02,1.960000000000000000e+02,1.970000000000000000e+02,1.970000000000000000e+02,1.970000000000000000e+02,1.970000000000000000e+02,1.970000000000000000e+02,1.980000000000000000e+02,1.970000000000000000e+02,1.960000000000000000e+02,1.980000000000000000e+02,1.960000000000000000e+02,1.960000000000000000e+02,1.930000000000000000e+02,1.970000000000000000e+02,1.970000000000000000e+02,1.970000000000000000e+02,1.970000000000000000e+02,1.970000000000000000e+02,1.940000000000000000e+02,1.940000000000000000e+02),
(5.900000000000000000e+01,5.100000000000000000e+01,7.600000000000000000e+01,9.500000000000000000e+01,8.800000000000000000e+01,6.600000000000000000e+01,6.100000000000000000e+01,6.700000000000000000e+01,5.800000000000000000e+01,1.130000000000000000e+02,1.210000000000000000e+02,9.900000000000000000e+01,8.800000000000000000e+01,8.200000000000000000e+01,1.260000000000000000e+02,1.490000000000000000e+02,8.400000000000000000e+01,1.800000000000000000e+01,1.700000000000000000e+01,3.300000000000000000e+01,4.500000000000000000e+01,6.700000000000000000e+01,9.200000000000000000e+01,1.180000000000000000e+02,1.150000000000000000e+02,1.220000000000000000e+02,1.040000000000000000e+02,8.400000000000000000e+01,9.500000000000000000e+01,1.370000000000000000e+02,1.510000000000000000e+02,1.570000000000000000e+02,1.670000000000000000e+02,1.870000000000000000e+02,1.990000000000000000e+02,2.020000000000000000e+02,2.080000000000000000e+02,1.940000000000000000e+02,1.610000000000000000e+02,1.650000000000000000e+02,1.860000000000000000e+02,1.960000000000000000e+02,1.920000000000000000e+02,1.840000000000000000e+02,1.560000000000000000e+02,1.410000000000000000e+02,9.900000000000000000e+01,6.900000000000000000e+01,6.000000000000000000e+01,3.400000000000000000e+01,9.700000000000000000e+01,1.190000000000000000e+02,1.180000000000000000e+02,1.480000000000000000e+02,1.750000000000000000e+02,1.790000000000000000e+02,1.820000000000000000e+02,1.650000000000000000e+02,1.940000000000000000e+02,1.830000000000000000e+02,1.880000000000000000e+02,1.950000000000000000e+02,1.840000000000000000e+02,1.990000000000000000e+02,1.910000000000000000e+02,2.090000000000000000e+02,2.090000000000000000e+02,2.110000000000000000e+02,2.090000000000000000e+02,2.080000000000000000e+02,2.030000000000000000e+02,2.070000000000000000e+02,2.090000000000000000e+02,2.090000000000000000e+02,2.110000000000000000e+02,2.070000000000000000e+02,2.080000000000000000e+02,2.070000000000000000e+02,2.100000000000000000e+02,2.030000000000000000e+02,2.090000000000000000e+02,1.920000000000000000e+02,2.020000000000000000e+02,1.700000000000000000e+02,1.570000000000000000e+02,6.100000000000000000e+01,3.900000000000000000e+01,3.700000000000000000e+01,2.100000000000000000e+01,2.400000000000000000e+01,6.700000000000000000e+01,6.300000000000000000e+01,8.700000000000000000e+01,1.280000000000000000e+02,1.100000000000000000e+02,1.020000000000000000e+02,6.700000000000000000e+01,7.400000000000000000e+01,1.310000000000000000e+02,4.200000000000000000e+01,2.800000000000000000e+01,6.200000000000000000e+01,6.400000000000000000e+01,1.320000000000000000e+02,1.750000000000000000e+02,1.960000000000000000e+02,1.980000000000000000e+02,1.980000000000000000e+02,1.970000000000000000e+02,2.020000000000000000e+02,2.030000000000000000e+02,2.030000000000000000e+02,2.030000000000000000e+02,2.030000000000000000e+02,2.020000000000000000e+02,2.040000000000000000e+02,2.010000000000000000e+02,2.020000000000000000e+02,2.020000000000000000e+02,2.020000000000000000e+02,1.980000000000000000e+02,2.000000000000000000e+02,2.010000000000000000e+02,2.020000000000000000e+02,2.000000000000000000e+02,2.000000000000000000e+02,2.000000000000000000e+02,2.000000000000000000e+02),
(6.600000000000000000e+01,5.100000000000000000e+01,8.300000000000000000e+01,1.210000000000000000e+02,9.700000000000000000e+01,5.500000000000000000e+01,6.600000000000000000e+01,6.700000000000000000e+01,7.100000000000000000e+01,7.500000000000000000e+01,1.200000000000000000e+02,1.130000000000000000e+02,8.200000000000000000e+01,1.430000000000000000e+02,1.260000000000000000e+02,8.100000000000000000e+01,1.000000000000000000e+02,3.600000000000000000e+01,1.500000000000000000e+01,4.000000000000000000e+01,6.100000000000000000e+01,6.500000000000000000e+01,6.600000000000000000e+01,6.000000000000000000e+01,9.100000000000000000e+01,1.150000000000000000e+02,1.480000000000000000e+02,1.400000000000000000e+02,1.240000000000000000e+02,1.020000000000000000e+02,1.450000000000000000e+02,1.550000000000000000e+02,1.820000000000000000e+02,1.770000000000000000e+02,1.920000000000000000e+02,1.980000000000000000e+02,1.840000000000000000e+02,1.980000000000000000e+02,1.900000000000000000e+02,2.000000000000000000e+02,1.990000000000000000e+02,2.070000000000000000e+02,2.020000000000000000e+02,1.820000000000000000e+02,1.670000000000000000e+02,1.580000000000000000e+02,1.290000000000000000e+02,1.270000000000000000e+02,7.500000000000000000e+01,7.500000000000000000e+01,8.100000000000000000e+01,1.030000000000000000e+02,1.130000000000000000e+02,1.540000000000000000e+02,1.330000000000000000e+02,1.890000000000000000e+02,1.870000000000000000e+02,1.820000000000000000e+02,1.820000000000000000e+02,1.630000000000000000e+02,1.840000000000000000e+02,1.870000000000000000e+02,1.920000000000000000e+02,1.790000000000000000e+02,1.820000000000000000e+02,1.960000000000000000e+02,2.020000000000000000e+02,2.070000000000000000e+02,1.990000000000000000e+02,1.990000000000000000e+02,2.000000000000000000e+02,2.050000000000000000e+02,2.090000000000000000e+02,2.080000000000000000e+02,2.100000000000000000e+02,1.980000000000000000e+02,2.040000000000000000e+02,2.020000000000000000e+02,2.100000000000000000e+02,1.840000000000000000e+02,2.070000000000000000e+02,2.020000000000000000e+02,1.300000000000000000e+02,1.020000000000000000e+02,5.100000000000000000e+01,2.400000000000000000e+01,2.400000000000000000e+01,9.000000000000000000e+00,2.500000000000000000e+01,4.000000000000000000e+01,9.300000000000000000e+01,8.600000000000000000e+01,8.700000000000000000e+01,1.050000000000000000e+02,1.030000000000000000e+02,7.800000000000000000e+01,6.700000000000000000e+01,3.000000000000000000e+01,4.000000000000000000e+01,7.400000000000000000e+01,4.300000000000000000e+01,6.700000000000000000e+01,1.020000000000000000e+02,9.600000000000000000e+01,1.600000000000000000e+02,1.860000000000000000e+02,1.950000000000000000e+02,2.010000000000000000e+02,2.050000000000000000e+02,2.030000000000000000e+02,2.050000000000000000e+02,2.060000000000000000e+02,2.060000000000000000e+02,2.060000000000000000e+02,2.050000000000000000e+02,2.050000000000000000e+02,2.050000000000000000e+02,2.050000000000000000e+02,2.050000000000000000e+02,2.040000000000000000e+02,2.030000000000000000e+02,2.020000000000000000e+02,2.050000000000000000e+02,2.050000000000000000e+02,2.050000000000000000e+02,2.040000000000000000e+02,2.030000000000000000e+02,2.000000000000000000e+02),
(5.100000000000000000e+01,5.200000000000000000e+01,1.070000000000000000e+02,1.350000000000000000e+02,1.080000000000000000e+02,7.400000000000000000e+01,4.700000000000000000e+01,3.200000000000000000e+01,4.600000000000000000e+01,4.400000000000000000e+01,5.900000000000000000e+01,6.200000000000000000e+01,6.900000000000000000e+01,1.100000000000000000e+02,1.230000000000000000e+02,9.600000000000000000e+01,7.500000000000000000e+01,3.600000000000000000e+01,1.500000000000000000e+01,1.100000000000000000e+01,1.700000000000000000e+01,5.500000000000000000e+01,1.400000000000000000e+01,3.000000000000000000e+01,1.160000000000000000e+02,1.440000000000000000e+02,1.580000000000000000e+02,1.430000000000000000e+02,1.270000000000000000e+02,1.080000000000000000e+02,1.060000000000000000e+02,1.150000000000000000e+02,1.100000000000000000e+02,1.250000000000000000e+02,1.750000000000000000e+02,1.760000000000000000e+02,1.970000000000000000e+02,1.710000000000000000e+02,1.970000000000000000e+02,1.870000000000000000e+02,2.020000000000000000e+02,1.890000000000000000e+02,1.720000000000000000e+02,1.560000000000000000e+02,1.680000000000000000e+02,1.980000000000000000e+02,1.860000000000000000e+02,1.530000000000000000e+02,1.350000000000000000e+02,1.380000000000000000e+02,9.100000000000000000e+01,1.070000000000000000e+02,1.290000000000000000e+02,1.360000000000000000e+02,1.040000000000000000e+02,1.830000000000000000e+02,1.270000000000000000e+02,1.710000000000000000e+02,1.470000000000000000e+02,1.320000000000000000e+02,1.590000000000000000e+02,1.660000000000000000e+02,1.740000000000000000e+02,1.670000000000000000e+02,1.660000000000000000e+02,1.810000000000000000e+02,1.780000000000000000e+02,1.910000000000000000e+02,1.930000000000000000e+02,1.930000000000000000e+02,1.970000000000000000e+02,2.050000000000000000e+02,2.030000000000000000e+02,2.010000000000000000e+02,2.070000000000000000e+02,1.930000000000000000e+02,1.890000000000000000e+02,1.970000000000000000e+02,1.840000000000000000e+02,1.840000000000000000e+02,1.720000000000000000e+02,1.480000000000000000e+02,9.100000000000000000e+01,2.500000000000000000e+01,1.700000000000000000e+01,1.400000000000000000e+01,3.900000000000000000e+01,1.000000000000000000e+01,2.600000000000000000e+01,3.700000000000000000e+01,8.500000000000000000e+01,7.900000000000000000e+01,9.400000000000000000e+01,1.000000000000000000e+02,1.400000000000000000e+02,1.030000000000000000e+02,3.100000000000000000e+01,1.500000000000000000e+01,8.000000000000000000e+00,7.000000000000000000e+01,7.900000000000000000e+01,7.200000000000000000e+01,8.500000000000000000e+01,1.050000000000000000e+02,1.590000000000000000e+02,1.900000000000000000e+02,1.960000000000000000e+02,1.960000000000000000e+02,1.990000000000000000e+02,1.970000000000000000e+02,1.950000000000000000e+02,1.980000000000000000e+02,1.970000000000000000e+02,1.970000000000000000e+02,1.980000000000000000e+02,1.980000000000000000e+02,1.970000000000000000e+02,1.970000000000000000e+02,1.960000000000000000e+02,1.950000000000000000e+02,1.960000000000000000e+02,1.910000000000000000e+02,1.950000000000000000e+02,1.950000000000000000e+02,1.940000000000000000e+02,1.940000000000000000e+02,1.940000000000000000e+02,1.910000000000000000e+02),
(4.400000000000000000e+01,8.100000000000000000e+01,1.260000000000000000e+02,1.260000000000000000e+02,1.210000000000000000e+02,8.100000000000000000e+01,3.900000000000000000e+01,4.800000000000000000e+01,4.900000000000000000e+01,6.600000000000000000e+01,6.700000000000000000e+01,7.000000000000000000e+01,1.020000000000000000e+02,9.600000000000000000e+01,1.280000000000000000e+02,8.600000000000000000e+01,5.400000000000000000e+01,2.900000000000000000e+01,1.100000000000000000e+01,1.000000000000000000e+01,5.400000000000000000e+01,1.600000000000000000e+01,4.200000000000000000e+01,9.000000000000000000e+01,1.490000000000000000e+02,1.500000000000000000e+02,1.430000000000000000e+02,1.740000000000000000e+02,1.420000000000000000e+02,1.050000000000000000e+02,9.500000000000000000e+01,8.100000000000000000e+01,9.300000000000000000e+01,1.500000000000000000e+02,1.490000000000000000e+02,1.590000000000000000e+02,1.500000000000000000e+02,1.780000000000000000e+02,1.760000000000000000e+02,1.590000000000000000e+02,1.560000000000000000e+02,1.680000000000000000e+02,1.410000000000000000e+02,1.880000000000000000e+02,1.970000000000000000e+02,1.590000000000000000e+02,1.260000000000000000e+02,1.400000000000000000e+02,1.660000000000000000e+02,1.710000000000000000e+02,1.280000000000000000e+02,1.440000000000000000e+02,1.650000000000000000e+02,1.200000000000000000e+02,1.150000000000000000e+02,1.540000000000000000e+02,1.560000000000000000e+02,1.600000000000000000e+02,1.450000000000000000e+02,1.350000000000000000e+02,1.580000000000000000e+02,1.620000000000000000e+02,1.650000000000000000e+02,1.740000000000000000e+02,1.580000000000000000e+02,1.670000000000000000e+02,1.620000000000000000e+02,1.930000000000000000e+02,1.730000000000000000e+02,1.950000000000000000e+02,1.900000000000000000e+02,1.870000000000000000e+02,1.900000000000000000e+02,1.620000000000000000e+02,1.830000000000000000e+02,1.820000000000000000e+02,1.720000000000000000e+02,1.960000000000000000e+02,1.590000000000000000e+02,1.240000000000000000e+02,7.000000000000000000e+01,9.500000000000000000e+01,1.350000000000000000e+02,2.200000000000000000e+01,1.500000000000000000e+01,1.900000000000000000e+01,3.700000000000000000e+01,2.300000000000000000e+01,2.400000000000000000e+01,2.700000000000000000e+01,7.500000000000000000e+01,6.400000000000000000e+01,4.400000000000000000e+01,4.300000000000000000e+01,4.300000000000000000e+01,8.800000000000000000e+01,1.700000000000000000e+01,1.200000000000000000e+01,1.900000000000000000e+01,3.700000000000000000e+01,8.800000000000000000e+01,5.600000000000000000e+01,6.500000000000000000e+01,9.600000000000000000e+01,1.280000000000000000e+02,1.650000000000000000e+02,1.860000000000000000e+02,1.860000000000000000e+02,1.890000000000000000e+02,1.940000000000000000e+02,1.850000000000000000e+02,1.820000000000000000e+02,1.850000000000000000e+02,1.830000000000000000e+02,1.860000000000000000e+02,1.850000000000000000e+02,1.890000000000000000e+02,1.820000000000000000e+02,1.880000000000000000e+02,1.820000000000000000e+02,1.820000000000000000e+02,1.830000000000000000e+02,1.840000000000000000e+02,1.840000000000000000e+02,1.810000000000000000e+02,1.830000000000000000e+02,1.820000000000000000e+02,1.810000000000000000e+02),
(6.500000000000000000e+01,8.900000000000000000e+01,9.400000000000000000e+01,1.230000000000000000e+02,1.400000000000000000e+02,7.700000000000000000e+01,3.700000000000000000e+01,5.200000000000000000e+01,5.900000000000000000e+01,5.700000000000000000e+01,6.400000000000000000e+01,8.000000000000000000e+01,9.200000000000000000e+01,1.110000000000000000e+02,1.630000000000000000e+02,1.570000000000000000e+02,8.600000000000000000e+01,5.900000000000000000e+01,2.000000000000000000e+01,3.100000000000000000e+01,5.000000000000000000e+00,2.000000000000000000e+00,5.000000000000000000e+00,2.800000000000000000e+01,3.100000000000000000e+01,5.600000000000000000e+01,8.100000000000000000e+01,9.500000000000000000e+01,1.130000000000000000e+02,1.390000000000000000e+02,1.100000000000000000e+02,7.400000000000000000e+01,1.260000000000000000e+02,9.300000000000000000e+01,1.210000000000000000e+02,1.410000000000000000e+02,1.620000000000000000e+02,1.710000000000000000e+02,1.540000000000000000e+02,1.420000000000000000e+02,1.670000000000000000e+02,1.620000000000000000e+02,1.730000000000000000e+02,1.650000000000000000e+02,1.130000000000000000e+02,1.230000000000000000e+02,1.410000000000000000e+02,1.750000000000000000e+02,1.600000000000000000e+02,1.500000000000000000e+02,1.920000000000000000e+02,1.900000000000000000e+02,1.690000000000000000e+02,7.900000000000000000e+01,8.300000000000000000e+01,1.370000000000000000e+02,1.530000000000000000e+02,1.010000000000000000e+02,1.600000000000000000e+02,1.540000000000000000e+02,1.460000000000000000e+02,1.600000000000000000e+02,1.540000000000000000e+02,1.560000000000000000e+02,1.480000000000000000e+02,1.370000000000000000e+02,1.500000000000000000e+02,1.930000000000000000e+02,1.630000000000000000e+02,1.760000000000000000e+02,1.720000000000000000e+02,1.640000000000000000e+02,1.490000000000000000e+02,1.410000000000000000e+02,1.380000000000000000e+02,1.380000000000000000e+02,1.480000000000000000e+02,1.390000000000000000e+02,1.490000000000000000e+02,6.500000000000000000e+01,4.300000000000000000e+01,2.800000000000000000e+01,9.500000000000000000e+01,1.600000000000000000e+01,9.000000000000000000e+00,1.600000000000000000e+01,1.400000000000000000e+01,2.200000000000000000e+01,4.300000000000000000e+01,3.500000000000000000e+01,4.100000000000000000e+01,3.800000000000000000e+01,3.100000000000000000e+01,3.000000000000000000e+01,1.000000000000000000e+01,5.600000000000000000e+01,1.700000000000000000e+01,2.100000000000000000e+01,4.000000000000000000e+01,5.200000000000000000e+01,6.600000000000000000e+01,8.000000000000000000e+01,8.500000000000000000e+01,1.000000000000000000e+02,1.130000000000000000e+02,1.270000000000000000e+02,1.500000000000000000e+02,1.730000000000000000e+02,1.640000000000000000e+02,1.710000000000000000e+02,1.700000000000000000e+02,1.650000000000000000e+02,1.640000000000000000e+02,1.650000000000000000e+02,1.660000000000000000e+02,1.640000000000000000e+02,1.640000000000000000e+02,1.650000000000000000e+02,1.660000000000000000e+02,1.630000000000000000e+02,1.640000000000000000e+02,1.640000000000000000e+02,1.640000000000000000e+02,1.640000000000000000e+02,1.610000000000000000e+02,1.590000000000000000e+02,1.600000000000000000e+02,1.610000000000000000e+02),
(5.400000000000000000e+01,9.800000000000000000e+01,1.250000000000000000e+02,1.150000000000000000e+02,1.150000000000000000e+02,7.600000000000000000e+01,3.500000000000000000e+01,3.800000000000000000e+01,5.100000000000000000e+01,6.400000000000000000e+01,6.500000000000000000e+01,8.000000000000000000e+01,1.040000000000000000e+02,1.620000000000000000e+02,1.330000000000000000e+02,1.340000000000000000e+02,1.010000000000000000e+02,6.100000000000000000e+01,2.700000000000000000e+01,4.700000000000000000e+01,1.500000000000000000e+01,1.000000000000000000e+01,1.600000000000000000e+01,1.300000000000000000e+01,4.000000000000000000e+01,7.500000000000000000e+01,1.180000000000000000e+02,1.480000000000000000e+02,1.510000000000000000e+02,1.400000000000000000e+02,1.360000000000000000e+02,1.590000000000000000e+02,1.090000000000000000e+02,1.240000000000000000e+02,1.290000000000000000e+02,1.290000000000000000e+02,1.560000000000000000e+02,1.340000000000000000e+02,1.390000000000000000e+02,1.570000000000000000e+02,1.580000000000000000e+02,1.850000000000000000e+02,1.540000000000000000e+02,1.330000000000000000e+02,1.460000000000000000e+02,1.710000000000000000e+02,1.480000000000000000e+02,1.140000000000000000e+02,1.850000000000000000e+02,1.900000000000000000e+02,1.380000000000000000e+02,1.870000000000000000e+02,1.280000000000000000e+02,1.030000000000000000e+02,8.500000000000000000e+01,1.180000000000000000e+02,1.220000000000000000e+02,8.300000000000000000e+01,1.470000000000000000e+02,1.490000000000000000e+02,1.380000000000000000e+02,1.600000000000000000e+02,1.310000000000000000e+02,1.560000000000000000e+02,1.340000000000000000e+02,1.290000000000000000e+02,1.430000000000000000e+02,1.490000000000000000e+02,1.460000000000000000e+02,1.510000000000000000e+02,1.470000000000000000e+02,1.360000000000000000e+02,1.180000000000000000e+02,9.400000000000000000e+01,9.100000000000000000e+01,7.900000000000000000e+01,9.900000000000000000e+01,4.400000000000000000e+01,7.300000000000000000e+01,4.200000000000000000e+01,1.900000000000000000e+01,2.800000000000000000e+01,1.400000000000000000e+01,1.320000000000000000e+02,2.500000000000000000e+01,2.600000000000000000e+01,1.500000000000000000e+01,1.700000000000000000e+01,3.300000000000000000e+01,4.100000000000000000e+01,2.800000000000000000e+01,1.300000000000000000e+01,6.000000000000000000e+00,6.000000000000000000e+00,1.000000000000000000e+01,4.000000000000000000e+00,3.000000000000000000e+01,3.700000000000000000e+01,5.700000000000000000e+01,7.700000000000000000e+01,8.500000000000000000e+01,1.280000000000000000e+02,1.090000000000000000e+02,8.200000000000000000e+01,7.900000000000000000e+01,7.600000000000000000e+01,9.300000000000000000e+01,1.210000000000000000e+02,1.440000000000000000e+02,1.350000000000000000e+02,1.590000000000000000e+02,1.330000000000000000e+02,1.260000000000000000e+02,1.290000000000000000e+02,1.260000000000000000e+02,1.270000000000000000e+02,1.280000000000000000e+02,1.250000000000000000e+02,1.350000000000000000e+02,1.260000000000000000e+02,1.270000000000000000e+02,1.220000000000000000e+02,1.200000000000000000e+02,1.260000000000000000e+02,1.250000000000000000e+02,1.250000000000000000e+02,1.240000000000000000e+02,1.160000000000000000e+02),
(6.700000000000000000e+01,1.510000000000000000e+02,1.490000000000000000e+02,1.060000000000000000e+02,8.300000000000000000e+01,6.300000000000000000e+01,3.900000000000000000e+01,5.200000000000000000e+01,5.100000000000000000e+01,5.200000000000000000e+01,1.180000000000000000e+02,1.360000000000000000e+02,1.210000000000000000e+02,1.210000000000000000e+02,1.690000000000000000e+02,1.860000000000000000e+02,1.600000000000000000e+02,1.200000000000000000e+02,7.100000000000000000e+01,2.000000000000000000e+01,1.100000000000000000e+01,8.000000000000000000e+00,1.200000000000000000e+01,5.200000000000000000e+01,2.800000000000000000e+01,4.000000000000000000e+01,7.800000000000000000e+01,9.600000000000000000e+01,9.000000000000000000e+01,9.000000000000000000e+01,1.270000000000000000e+02,1.590000000000000000e+02,1.710000000000000000e+02,1.590000000000000000e+02,1.590000000000000000e+02,1.230000000000000000e+02,1.100000000000000000e+02,9.900000000000000000e+01,1.340000000000000000e+02,1.530000000000000000e+02,1.240000000000000000e+02,1.690000000000000000e+02,1.840000000000000000e+02,1.700000000000000000e+02,1.800000000000000000e+02,1.760000000000000000e+02,1.550000000000000000e+02,1.620000000000000000e+02,1.720000000000000000e+02,1.730000000000000000e+02,1.800000000000000000e+02,1.400000000000000000e+02,1.740000000000000000e+02,1.280000000000000000e+02,1.410000000000000000e+02,1.080000000000000000e+02,9.500000000000000000e+01,6.500000000000000000e+01,1.230000000000000000e+02,1.380000000000000000e+02,1.150000000000000000e+02,1.270000000000000000e+02,1.250000000000000000e+02,1.260000000000000000e+02,1.210000000000000000e+02,1.100000000000000000e+02,1.180000000000000000e+02,1.220000000000000000e+02,1.310000000000000000e+02,1.020000000000000000e+02,9.400000000000000000e+01,8.500000000000000000e+01,9.000000000000000000e+01,4.400000000000000000e+01,4.800000000000000000e+01,3.500000000000000000e+01,3.400000000000000000e+01,4.100000000000000000e+01,2.300000000000000000e+01,2.800000000000000000e+01,1.900000000000000000e+01,5.100000000000000000e+01,2.400000000000000000e+01,2.100000000000000000e+01,8.900000000000000000e+01,2.200000000000000000e+01,1.500000000000000000e+01,1.800000000000000000e+01,9.000000000000000000e+00,2.000000000000000000e+00,4.000000000000000000e+00,6.000000000000000000e+00,2.000000000000000000e+00,2.000000000000000000e+00,5.000000000000000000e+00,4.000000000000000000e+00,6.300000000000000000e+01,3.700000000000000000e+01,5.400000000000000000e+01,6.200000000000000000e+01,7.300000000000000000e+01,1.080000000000000000e+02,8.800000000000000000e+01,7.400000000000000000e+01,5.700000000000000000e+01,4.900000000000000000e+01,5.400000000000000000e+01,7.200000000000000000e+01,8.200000000000000000e+01,8.800000000000000000e+01,9.000000000000000000e+01,1.210000000000000000e+02,7.400000000000000000e+01,7.500000000000000000e+01,7.800000000000000000e+01,7.800000000000000000e+01,7.500000000000000000e+01,7.500000000000000000e+01,7.300000000000000000e+01,7.900000000000000000e+01,7.000000000000000000e+01,7.300000000000000000e+01,7.500000000000000000e+01,7.500000000000000000e+01,7.700000000000000000e+01,7.400000000000000000e+01,7.200000000000000000e+01,7.200000000000000000e+01),
(9.900000000000000000e+01,1.630000000000000000e+02,1.560000000000000000e+02,1.360000000000000000e+02,8.800000000000000000e+01,7.900000000000000000e+01,5.000000000000000000e+01,2.800000000000000000e+01,4.500000000000000000e+01,6.900000000000000000e+01,7.500000000000000000e+01,1.230000000000000000e+02,1.120000000000000000e+02,1.150000000000000000e+02,1.400000000000000000e+02,1.630000000000000000e+02,1.440000000000000000e+02,1.130000000000000000e+02,7.900000000000000000e+01,3.100000000000000000e+01,1.300000000000000000e+01,1.500000000000000000e+01,1.300000000000000000e+01,1.000000000000000000e+01,2.800000000000000000e+01,3.700000000000000000e+01,3.100000000000000000e+01,6.700000000000000000e+01,9.500000000000000000e+01,1.300000000000000000e+02,1.860000000000000000e+02,1.710000000000000000e+02,1.590000000000000000e+02,1.640000000000000000e+02,1.340000000000000000e+02,1.160000000000000000e+02,1.590000000000000000e+02,1.720000000000000000e+02,1.550000000000000000e+02,1.550000000000000000e+02,1.530000000000000000e+02,1.570000000000000000e+02,1.650000000000000000e+02,1.910000000000000000e+02,1.740000000000000000e+02,1.590000000000000000e+02,1.450000000000000000e+02,1.590000000000000000e+02,1.840000000000000000e+02,1.750000000000000000e+02,1.610000000000000000e+02,1.690000000000000000e+02,1.700000000000000000e+02,1.810000000000000000e+02,1.610000000000000000e+02,1.700000000000000000e+02,9.200000000000000000e+01,5.600000000000000000e+01,1.510000000000000000e+02,1.050000000000000000e+02,8.800000000000000000e+01,9.800000000000000000e+01,8.900000000000000000e+01,9.600000000000000000e+01,8.600000000000000000e+01,6.200000000000000000e+01,9.000000000000000000e+01,7.000000000000000000e+01,7.700000000000000000e+01,3.700000000000000000e+01,4.800000000000000000e+01,2.200000000000000000e+01,2.400000000000000000e+01,4.000000000000000000e+01,1.900000000000000000e+01,3.000000000000000000e+01,1.900000000000000000e+01,5.700000000000000000e+01,2.100000000000000000e+01,2.500000000000000000e+01,1.500000000000000000e+01,1.600000000000000000e+01,5.200000000000000000e+01,7.000000000000000000e+00,5.000000000000000000e+00,1.600000000000000000e+01,3.000000000000000000e+00,1.000000000000000000e+00,2.000000000000000000e+00,2.000000000000000000e+00,2.000000000000000000e+00,2.000000000000000000e+00,3.000000000000000000e+00,5.000000000000000000e+00,5.000000000000000000e+00,9.000000000000000000e+00,5.100000000000000000e+01,7.800000000000000000e+01,8.300000000000000000e+01,6.300000000000000000e+01,5.600000000000000000e+01,6.200000000000000000e+01,7.300000000000000000e+01,4.500000000000000000e+01,4.400000000000000000e+01,2.800000000000000000e+01,2.500000000000000000e+01,2.800000000000000000e+01,2.800000000000000000e+01,4.700000000000000000e+01,2.700000000000000000e+01,3.900000000000000000e+01,6.200000000000000000e+01,2.600000000000000000e+01,2.700000000000000000e+01,2.700000000000000000e+01,2.600000000000000000e+01,2.900000000000000000e+01,2.800000000000000000e+01,2.800000000000000000e+01,2.500000000000000000e+01,2.500000000000000000e+01,2.600000000000000000e+01,2.600000000000000000e+01,2.600000000000000000e+01,2.800000000000000000e+01,2.900000000000000000e+01,2.600000000000000000e+01),
(1.030000000000000000e+02,1.700000000000000000e+02,1.730000000000000000e+02,1.400000000000000000e+02,1.210000000000000000e+02,9.300000000000000000e+01,6.200000000000000000e+01,5.500000000000000000e+01,4.400000000000000000e+01,4.900000000000000000e+01,4.800000000000000000e+01,8.500000000000000000e+01,1.360000000000000000e+02,1.460000000000000000e+02,1.210000000000000000e+02,1.280000000000000000e+02,1.470000000000000000e+02,1.300000000000000000e+02,7.200000000000000000e+01,2.700000000000000000e+01,1.900000000000000000e+01,1.200000000000000000e+01,1.200000000000000000e+01,1.300000000000000000e+01,1.100000000000000000e+01,1.600000000000000000e+01,3.100000000000000000e+01,5.300000000000000000e+01,4.400000000000000000e+01,1.120000000000000000e+02,1.170000000000000000e+02,1.330000000000000000e+02,1.630000000000000000e+02,1.590000000000000000e+02,1.720000000000000000e+02,1.730000000000000000e+02,1.450000000000000000e+02,1.490000000000000000e+02,1.540000000000000000e+02,1.450000000000000000e+02,1.410000000000000000e+02,1.500000000000000000e+02,1.670000000000000000e+02,1.620000000000000000e+02,1.500000000000000000e+02,1.660000000000000000e+02,1.700000000000000000e+02,1.730000000000000000e+02,1.610000000000000000e+02,1.500000000000000000e+02,1.390000000000000000e+02,1.700000000000000000e+02,1.740000000000000000e+02,1.820000000000000000e+02,1.680000000000000000e+02,1.880000000000000000e+02,1.090000000000000000e+02,7.000000000000000000e+01,1.510000000000000000e+02,1.040000000000000000e+02,7.600000000000000000e+01,7.800000000000000000e+01,9.700000000000000000e+01,8.500000000000000000e+01,6.900000000000000000e+01,4.300000000000000000e+01,5.900000000000000000e+01,3.300000000000000000e+01,4.000000000000000000e+01,2.000000000000000000e+01,2.800000000000000000e+01,9.000000000000000000e+00,1.400000000000000000e+01,2.200000000000000000e+01,3.500000000000000000e+01,2.300000000000000000e+01,2.500000000000000000e+01,2.400000000000000000e+01,1.900000000000000000e+01,7.000000000000000000e+00,6.000000000000000000e+00,5.000000000000000000e+00,1.000000000000000000e+01,2.600000000000000000e+01,3.000000000000000000e+00,3.000000000000000000e+00,3.000000000000000000e+00,1.000000000000000000e+00,2.000000000000000000e+00,2.000000000000000000e+00,6.000000000000000000e+00,2.000000000000000000e+00,6.000000000000000000e+00,7.000000000000000000e+00,9.000000000000000000e+00,2.200000000000000000e+01,8.200000000000000000e+01,1.140000000000000000e+02,1.230000000000000000e+02,1.180000000000000000e+02,6.900000000000000000e+01,4.200000000000000000e+01,8.000000000000000000e+01,4.400000000000000000e+01,3.400000000000000000e+01,1.100000000000000000e+01,6.000000000000000000e+00,6.000000000000000000e+00,3.000000000000000000e+00,6.000000000000000000e+00,2.400000000000000000e+01,1.200000000000000000e+01,3.300000000000000000e+01,1.300000000000000000e+01,5.000000000000000000e+00,5.000000000000000000e+00,5.000000000000000000e+00,5.000000000000000000e+00,9.000000000000000000e+00,9.000000000000000000e+00,6.000000000000000000e+00,6.000000000000000000e+00,4.000000000000000000e+00,7.000000000000000000e+00,1.000000000000000000e+01,9.000000000000000000e+00,9.000000000000000000e+00,9.000000000000000000e+00),
(1.070000000000000000e+02,1.640000000000000000e+02,1.790000000000000000e+02,1.550000000000000000e+02,1.030000000000000000e+02,9.200000000000000000e+01,8.300000000000000000e+01,4.200000000000000000e+01,2.000000000000000000e+01,2.000000000000000000e+01,3.000000000000000000e+01,7.300000000000000000e+01,6.800000000000000000e+01,9.400000000000000000e+01,1.380000000000000000e+02,1.340000000000000000e+02,1.580000000000000000e+02,1.820000000000000000e+02,1.590000000000000000e+02,4.800000000000000000e+01,2.900000000000000000e+01,2.700000000000000000e+01,1.300000000000000000e+01,1.200000000000000000e+01,8.000000000000000000e+00,1.500000000000000000e+01,3.500000000000000000e+01,4.500000000000000000e+01,4.400000000000000000e+01,1.240000000000000000e+02,1.030000000000000000e+02,1.390000000000000000e+02,1.320000000000000000e+02,1.260000000000000000e+02,1.410000000000000000e+02,1.650000000000000000e+02,1.500000000000000000e+02,1.730000000000000000e+02,1.220000000000000000e+02,1.010000000000000000e+02,1.400000000000000000e+02,1.840000000000000000e+02,1.850000000000000000e+02,1.710000000000000000e+02,1.890000000000000000e+02,2.010000000000000000e+02,1.660000000000000000e+02,1.700000000000000000e+02,1.770000000000000000e+02,1.190000000000000000e+02,1.590000000000000000e+02,1.990000000000000000e+02,1.780000000000000000e+02,1.750000000000000000e+02,1.910000000000000000e+02,1.880000000000000000e+02,1.520000000000000000e+02,1.020000000000000000e+02,1.350000000000000000e+02,1.280000000000000000e+02,8.500000000000000000e+01,9.800000000000000000e+01,1.040000000000000000e+02,1.150000000000000000e+02,9.200000000000000000e+01,8.300000000000000000e+01,5.500000000000000000e+01,2.800000000000000000e+01,3.800000000000000000e+01,2.100000000000000000e+01,2.300000000000000000e+01,2.400000000000000000e+01,1.800000000000000000e+01,2.200000000000000000e+01,2.700000000000000000e+01,3.300000000000000000e+01,3.700000000000000000e+01,2.100000000000000000e+01,1.800000000000000000e+01,1.000000000000000000e+01,6.000000000000000000e+00,3.000000000000000000e+00,4.000000000000000000e+00,4.000000000000000000e+00,5.000000000000000000e+00,8.000000000000000000e+00,5.000000000000000000e+00,3.000000000000000000e+00,3.000000000000000000e+00,4.000000000000000000e+00,4.000000000000000000e+00,5.000000000000000000e+00,6.000000000000000000e+00,1.100000000000000000e+01,2.800000000000000000e+01,5.600000000000000000e+01,8.000000000000000000e+01,1.520000000000000000e+02,1.250000000000000000e+02,9.700000000000000000e+01,9.400000000000000000e+01,9.600000000000000000e+01,9.400000000000000000e+01,4.400000000000000000e+01,1.800000000000000000e+01,5.000000000000000000e+00,2.000000000000000000e+00,0.000000000000000000e+00,1.000000000000000000e+00,1.000000000000000000e+00,2.000000000000000000e+00,6.000000000000000000e+00,5.000000000000000000e+00,1.400000000000000000e+01,4.000000000000000000e+00,1.000000000000000000e+00,1.000000000000000000e+00,1.000000000000000000e+00,1.000000000000000000e+00,2.000000000000000000e+00,2.000000000000000000e+00,3.000000000000000000e+00,3.000000000000000000e+00,1.000000000000000000e+00,3.000000000000000000e+00,3.000000000000000000e+00,3.000000000000000000e+00,3.000000000000000000e+00),
(9.400000000000000000e+01,1.890000000000000000e+02,1.870000000000000000e+02,1.640000000000000000e+02,1.250000000000000000e+02,9.100000000000000000e+01,7.000000000000000000e+01,7.000000000000000000e+01,3.900000000000000000e+01,3.000000000000000000e+01,2.000000000000000000e+01,6.200000000000000000e+01,9.700000000000000000e+01,7.700000000000000000e+01,9.600000000000000000e+01,1.250000000000000000e+02,1.730000000000000000e+02,1.730000000000000000e+02,1.620000000000000000e+02,1.000000000000000000e+02,5.500000000000000000e+01,2.500000000000000000e+01,1.300000000000000000e+01,2.100000000000000000e+01,2.000000000000000000e+01,1.200000000000000000e+01,2.000000000000000000e+01,3.400000000000000000e+01,8.600000000000000000e+01,9.900000000000000000e+01,1.610000000000000000e+02,1.610000000000000000e+02,1.610000000000000000e+02,1.670000000000000000e+02,1.770000000000000000e+02,1.260000000000000000e+02,9.900000000000000000e+01,1.480000000000000000e+02,1.280000000000000000e+02,1.100000000000000000e+02,1.600000000000000000e+02,1.810000000000000000e+02,1.520000000000000000e+02,1.840000000000000000e+02,1.930000000000000000e+02,1.540000000000000000e+02,1.670000000000000000e+02,2.020000000000000000e+02,1.640000000000000000e+02,1.300000000000000000e+02,1.780000000000000000e+02,1.800000000000000000e+02,1.900000000000000000e+02,1.810000000000000000e+02,1.790000000000000000e+02,1.690000000000000000e+02,1.550000000000000000e+02,1.490000000000000000e+02,1.350000000000000000e+02,1.510000000000000000e+02,1.410000000000000000e+02,1.250000000000000000e+02,1.100000000000000000e+02,1.210000000000000000e+02,1.390000000000000000e+02,1.090000000000000000e+02,7.500000000000000000e+01,8.900000000000000000e+01,5.800000000000000000e+01,5.200000000000000000e+01,5.500000000000000000e+01,3.900000000000000000e+01,2.500000000000000000e+01,3.500000000000000000e+01,2.700000000000000000e+01,2.200000000000000000e+01,1.500000000000000000e+01,2.000000000000000000e+01,1.200000000000000000e+01,5.000000000000000000e+00,2.000000000000000000e+00,2.000000000000000000e+00,1.000000000000000000e+00,4.000000000000000000e+00,4.000000000000000000e+00,1.200000000000000000e+01,1.400000000000000000e+01,1.500000000000000000e+01,1.600000000000000000e+01,6.000000000000000000e+00,9.000000000000000000e+00,7.000000000000000000e+00,1.400000000000000000e+01,2.400000000000000000e+01,5.100000000000000000e+01,6.200000000000000000e+01,6.000000000000000000e+01,8.300000000000000000e+01,1.170000000000000000e+02,8.700000000000000000e+01,6.500000000000000000e+01,4.200000000000000000e+01,7.000000000000000000e+01,6.200000000000000000e+01,3.000000000000000000e+01,8.000000000000000000e+00,2.000000000000000000e+00,0.000000000000000000e+00,1.000000000000000000e+00,1.000000000000000000e+00,0.000000000000000000e+00,1.000000000000000000e+00,5.000000000000000000e+00,8.000000000000000000e+00,1.000000000000000000e+01,1.000000000000000000e+00,1.000000000000000000e+00,1.000000000000000000e+00,2.000000000000000000e+00,4.000000000000000000e+00,5.000000000000000000e+00,3.000000000000000000e+00,3.000000000000000000e+00,1.000000000000000000e+00,3.000000000000000000e+00,3.000000000000000000e+00,5.000000000000000000e+00,5.000000000000000000e+00),
(1.390000000000000000e+02,1.800000000000000000e+02,1.860000000000000000e+02,1.410000000000000000e+02,1.250000000000000000e+02,1.080000000000000000e+02,1.010000000000000000e+02,7.000000000000000000e+01,4.300000000000000000e+01,2.000000000000000000e+01,1.600000000000000000e+01,4.900000000000000000e+01,9.800000000000000000e+01,1.360000000000000000e+02,1.380000000000000000e+02,1.200000000000000000e+02,1.250000000000000000e+02,1.650000000000000000e+02,1.420000000000000000e+02,1.350000000000000000e+02,8.300000000000000000e+01,3.400000000000000000e+01,2.000000000000000000e+01,2.400000000000000000e+01,2.600000000000000000e+01,2.200000000000000000e+01,2.300000000000000000e+01,3.800000000000000000e+01,7.800000000000000000e+01,1.070000000000000000e+02,1.320000000000000000e+02,9.900000000000000000e+01,7.700000000000000000e+01,8.500000000000000000e+01,1.040000000000000000e+02,1.190000000000000000e+02,1.130000000000000000e+02,1.460000000000000000e+02,1.350000000000000000e+02,1.470000000000000000e+02,1.570000000000000000e+02,1.620000000000000000e+02,1.690000000000000000e+02,1.970000000000000000e+02,1.730000000000000000e+02,1.440000000000000000e+02,2.020000000000000000e+02,2.000000000000000000e+02,1.520000000000000000e+02,1.150000000000000000e+02,1.610000000000000000e+02,1.560000000000000000e+02,2.020000000000000000e+02,1.910000000000000000e+02,1.490000000000000000e+02,1.560000000000000000e+02,1.700000000000000000e+02,1.800000000000000000e+02,1.560000000000000000e+02,1.410000000000000000e+02,1.660000000000000000e+02,1.280000000000000000e+02,1.450000000000000000e+02,1.350000000000000000e+02,1.210000000000000000e+02,1.370000000000000000e+02,1.200000000000000000e+02,8.100000000000000000e+01,1.080000000000000000e+02,7.200000000000000000e+01,7.300000000000000000e+01,1.090000000000000000e+02,5.200000000000000000e+01,2.900000000000000000e+01,2.800000000000000000e+01,2.800000000000000000e+01,9.000000000000000000e+00,9.000000000000000000e+00,4.000000000000000000e+00,0.000000000000000000e+00,1.000000000000000000e+00,1.000000000000000000e+00,3.000000000000000000e+00,5.000000000000000000e+00,6.000000000000000000e+00,7.000000000000000000e+00,9.000000000000000000e+00,1.200000000000000000e+01,1.400000000000000000e+01,1.000000000000000000e+01,2.900000000000000000e+01,2.300000000000000000e+01,3.200000000000000000e+01,4.800000000000000000e+01,9.200000000000000000e+01,1.090000000000000000e+02,8.300000000000000000e+01,5.900000000000000000e+01,6.800000000000000000e+01,3.600000000000000000e+01,2.700000000000000000e+01,2.200000000000000000e+01,4.700000000000000000e+01,5.400000000000000000e+01,3.900000000000000000e+01,1.300000000000000000e+01,3.000000000000000000e+00,1.000000000000000000e+00,1.000000000000000000e+00,1.000000000000000000e+00,2.000000000000000000e+00,2.000000000000000000e+00,3.000000000000000000e+00,7.000000000000000000e+00,7.000000000000000000e+00,5.000000000000000000e+00,3.000000000000000000e+00,2.000000000000000000e+00,2.000000000000000000e+00,6.000000000000000000e+00,4.000000000000000000e+00,4.000000000000000000e+00,4.000000000000000000e+00,4.000000000000000000e+00,4.000000000000000000e+00,7.000000000000000000e+00,7.000000000000000000e+00,7.000000000000000000e+00),
(1.280000000000000000e+02,1.880000000000000000e+02,1.810000000000000000e+02,1.520000000000000000e+02,1.180000000000000000e+02,1.380000000000000000e+02,1.490000000000000000e+02,1.170000000000000000e+02,4.900000000000000000e+01,1.600000000000000000e+01,8.000000000000000000e+00,1.000000000000000000e+01,3.000000000000000000e+01,6.600000000000000000e+01,1.240000000000000000e+02,1.320000000000000000e+02,1.730000000000000000e+02,1.700000000000000000e+02,1.650000000000000000e+02,1.450000000000000000e+02,9.900000000000000000e+01,5.400000000000000000e+01,3.400000000000000000e+01,2.500000000000000000e+01,1.300000000000000000e+01,2.300000000000000000e+01,8.000000000000000000e+00,8.000000000000000000e+00,2.900000000000000000e+01,3.100000000000000000e+01,2.000000000000000000e+01,1.700000000000000000e+01,5.700000000000000000e+01,9.600000000000000000e+01,1.030000000000000000e+02,1.160000000000000000e+02,1.130000000000000000e+02,1.700000000000000000e+02,1.860000000000000000e+02,1.610000000000000000e+02,1.420000000000000000e+02,1.560000000000000000e+02,1.850000000000000000e+02,1.450000000000000000e+02,1.510000000000000000e+02,1.970000000000000000e+02,1.950000000000000000e+02,1.650000000000000000e+02,1.480000000000000000e+02,1.370000000000000000e+02,1.600000000000000000e+02,1.600000000000000000e+02,2.000000000000000000e+02,1.810000000000000000e+02,1.410000000000000000e+02,1.680000000000000000e+02,1.710000000000000000e+02,1.650000000000000000e+02,1.750000000000000000e+02,1.700000000000000000e+02,1.760000000000000000e+02,1.540000000000000000e+02,1.460000000000000000e+02,1.550000000000000000e+02,1.460000000000000000e+02,1.300000000000000000e+02,1.540000000000000000e+02,1.140000000000000000e+02,7.300000000000000000e+01,1.420000000000000000e+02,5.100000000000000000e+01,6.400000000000000000e+01,1.220000000000000000e+02,6.500000000000000000e+01,5.000000000000000000e+01,4.600000000000000000e+01,6.000000000000000000e+00,1.000000000000000000e+00,1.000000000000000000e+00,3.000000000000000000e+00,3.000000000000000000e+00,1.100000000000000000e+01,1.200000000000000000e+01,1.600000000000000000e+01,1.000000000000000000e+01,1.400000000000000000e+01,2.400000000000000000e+01,7.000000000000000000e+00,1.600000000000000000e+01,1.200000000000000000e+01,1.900000000000000000e+01,5.600000000000000000e+01,1.070000000000000000e+02,1.460000000000000000e+02,1.260000000000000000e+02,1.330000000000000000e+02,1.520000000000000000e+02,1.320000000000000000e+02,1.230000000000000000e+02,8.300000000000000000e+01,5.000000000000000000e+01,3.400000000000000000e+01,6.300000000000000000e+01,7.400000000000000000e+01,3.100000000000000000e+01,1.300000000000000000e+01,6.000000000000000000e+00,6.000000000000000000e+00,7.000000000000000000e+00,7.000000000000000000e+00,6.000000000000000000e+00,6.000000000000000000e+00,6.000000000000000000e+00,8.000000000000000000e+00,1.800000000000000000e+01,2.200000000000000000e+01,1.100000000000000000e+01,8.000000000000000000e+00,1.400000000000000000e+01,1.400000000000000000e+01,1.300000000000000000e+01,1.300000000000000000e+01,1.000000000000000000e+01,1.000000000000000000e+01,1.300000000000000000e+01,1.200000000000000000e+01,1.300000000000000000e+01,1.300000000000000000e+01),
(1.810000000000000000e+02,2.020000000000000000e+02,1.930000000000000000e+02,1.670000000000000000e+02,1.690000000000000000e+02,1.550000000000000000e+02,1.270000000000000000e+02,1.280000000000000000e+02,6.800000000000000000e+01,3.300000000000000000e+01,1.000000000000000000e+01,1.000000000000000000e+01,2.100000000000000000e+01,4.100000000000000000e+01,9.400000000000000000e+01,1.490000000000000000e+02,1.600000000000000000e+02,1.590000000000000000e+02,1.770000000000000000e+02,1.860000000000000000e+02,1.440000000000000000e+02,8.000000000000000000e+01,4.400000000000000000e+01,2.500000000000000000e+01,3.100000000000000000e+01,2.400000000000000000e+01,1.300000000000000000e+01,1.300000000000000000e+01,5.000000000000000000e+00,8.000000000000000000e+00,1.700000000000000000e+01,4.500000000000000000e+01,7.600000000000000000e+01,8.800000000000000000e+01,1.370000000000000000e+02,1.590000000000000000e+02,1.870000000000000000e+02,1.990000000000000000e+02,1.770000000000000000e+02,1.750000000000000000e+02,1.880000000000000000e+02,1.710000000000000000e+02,1.530000000000000000e+02,1.640000000000000000e+02,1.860000000000000000e+02,1.710000000000000000e+02,1.710000000000000000e+02,1.690000000000000000e+02,1.800000000000000000e+02,1.660000000000000000e+02,1.370000000000000000e+02,1.550000000000000000e+02,1.950000000000000000e+02,1.690000000000000000e+02,1.640000000000000000e+02,1.300000000000000000e+02,1.700000000000000000e+02,1.470000000000000000e+02,1.600000000000000000e+02,1.180000000000000000e+02,1.680000000000000000e+02,1.590000000000000000e+02,1.480000000000000000e+02,1.560000000000000000e+02,1.610000000000000000e+02,1.190000000000000000e+02,1.540000000000000000e+02,1.660000000000000000e+02,1.070000000000000000e+02,9.900000000000000000e+01,1.160000000000000000e+02,6.800000000000000000e+01,9.000000000000000000e+01,6.500000000000000000e+01,3.700000000000000000e+01,1.100000000000000000e+01,3.000000000000000000e+00,5.000000000000000000e+00,9.000000000000000000e+00,1.400000000000000000e+01,3.800000000000000000e+01,2.900000000000000000e+01,3.500000000000000000e+01,4.500000000000000000e+01,1.200000000000000000e+01,1.300000000000000000e+01,2.300000000000000000e+01,1.300000000000000000e+01,1.500000000000000000e+01,4.900000000000000000e+01,5.500000000000000000e+01,6.600000000000000000e+01,1.100000000000000000e+02,1.630000000000000000e+02,1.700000000000000000e+02,1.660000000000000000e+02,1.160000000000000000e+02,6.900000000000000000e+01,6.900000000000000000e+01,6.000000000000000000e+01,6.000000000000000000e+01,8.700000000000000000e+01,1.070000000000000000e+02,9.800000000000000000e+01,6.200000000000000000e+01,2.500000000000000000e+01,1.300000000000000000e+01,1.400000000000000000e+01,1.600000000000000000e+01,1.800000000000000000e+01,1.800000000000000000e+01,1.700000000000000000e+01,1.900000000000000000e+01,1.600000000000000000e+01,1.900000000000000000e+01,2.600000000000000000e+01,3.100000000000000000e+01,2.300000000000000000e+01,2.700000000000000000e+01,2.700000000000000000e+01,2.700000000000000000e+01,2.200000000000000000e+01,2.300000000000000000e+01,2.300000000000000000e+01,2.200000000000000000e+01,2.500000000000000000e+01,2.600000000000000000e+01,2.500000000000000000e+01),
(1.690000000000000000e+02,1.990000000000000000e+02,1.920000000000000000e+02,1.800000000000000000e+02,1.530000000000000000e+02,1.240000000000000000e+02,1.200000000000000000e+02,1.430000000000000000e+02,9.700000000000000000e+01,5.800000000000000000e+01,1.600000000000000000e+01,1.400000000000000000e+01,4.000000000000000000e+00,1.300000000000000000e+01,3.300000000000000000e+01,9.300000000000000000e+01,1.310000000000000000e+02,1.340000000000000000e+02,1.530000000000000000e+02,1.590000000000000000e+02,1.510000000000000000e+02,8.200000000000000000e+01,4.700000000000000000e+01,1.000000000000000000e+01,9.000000000000000000e+00,1.300000000000000000e+01,8.000000000000000000e+00,1.100000000000000000e+01,8.000000000000000000e+00,2.300000000000000000e+01,2.600000000000000000e+01,5.900000000000000000e+01,1.150000000000000000e+02,9.500000000000000000e+01,1.420000000000000000e+02,1.750000000000000000e+02,2.020000000000000000e+02,1.780000000000000000e+02,1.650000000000000000e+02,1.950000000000000000e+02,1.700000000000000000e+02,1.360000000000000000e+02,1.450000000000000000e+02,1.960000000000000000e+02,1.790000000000000000e+02,1.560000000000000000e+02,1.830000000000000000e+02,1.970000000000000000e+02,1.850000000000000000e+02,1.790000000000000000e+02,1.710000000000000000e+02,1.870000000000000000e+02,1.750000000000000000e+02,1.570000000000000000e+02,1.750000000000000000e+02,1.600000000000000000e+02,1.690000000000000000e+02,1.370000000000000000e+02,1.310000000000000000e+02,1.090000000000000000e+02,1.200000000000000000e+02,1.750000000000000000e+02,1.370000000000000000e+02,1.700000000000000000e+02,1.550000000000000000e+02,1.380000000000000000e+02,1.140000000000000000e+02,1.400000000000000000e+02,1.670000000000000000e+02,1.070000000000000000e+02,1.130000000000000000e+02,8.300000000000000000e+01,7.600000000000000000e+01,2.000000000000000000e+01,3.700000000000000000e+01,8.000000000000000000e+00,6.000000000000000000e+00,1.000000000000000000e+01,2.600000000000000000e+01,3.000000000000000000e+01,2.400000000000000000e+01,1.900000000000000000e+01,1.400000000000000000e+01,1.300000000000000000e+01,2.300000000000000000e+01,1.300000000000000000e+01,2.200000000000000000e+01,3.400000000000000000e+01,4.000000000000000000e+01,4.100000000000000000e+01,9.300000000000000000e+01,1.520000000000000000e+02,1.660000000000000000e+02,1.660000000000000000e+02,1.610000000000000000e+02,1.370000000000000000e+02,1.230000000000000000e+02,1.300000000000000000e+02,9.100000000000000000e+01,7.800000000000000000e+01,5.100000000000000000e+01,5.900000000000000000e+01,9.100000000000000000e+01,1.250000000000000000e+02,8.700000000000000000e+01,4.500000000000000000e+01,3.300000000000000000e+01,3.600000000000000000e+01,3.900000000000000000e+01,4.000000000000000000e+01,4.000000000000000000e+01,4.200000000000000000e+01,4.100000000000000000e+01,4.100000000000000000e+01,3.900000000000000000e+01,5.400000000000000000e+01,5.500000000000000000e+01,4.300000000000000000e+01,4.700000000000000000e+01,4.700000000000000000e+01,5.000000000000000000e+01,4.900000000000000000e+01,4.900000000000000000e+01,4.900000000000000000e+01,4.800000000000000000e+01,4.500000000000000000e+01,5.000000000000000000e+01,5.100000000000000000e+01),
(1.780000000000000000e+02,2.060000000000000000e+02,2.050000000000000000e+02,1.890000000000000000e+02,1.860000000000000000e+02,1.430000000000000000e+02,1.460000000000000000e+02,1.700000000000000000e+02,1.350000000000000000e+02,8.800000000000000000e+01,2.100000000000000000e+01,1.300000000000000000e+01,1.200000000000000000e+01,1.000000000000000000e+01,2.500000000000000000e+01,7.200000000000000000e+01,1.220000000000000000e+02,1.600000000000000000e+02,1.680000000000000000e+02,1.580000000000000000e+02,1.600000000000000000e+02,1.320000000000000000e+02,6.300000000000000000e+01,2.200000000000000000e+01,2.500000000000000000e+01,2.900000000000000000e+01,2.500000000000000000e+01,1.100000000000000000e+01,1.000000000000000000e+01,1.000000000000000000e+01,7.000000000000000000e+00,2.200000000000000000e+01,7.300000000000000000e+01,1.120000000000000000e+02,4.800000000000000000e+01,6.900000000000000000e+01,8.500000000000000000e+01,1.690000000000000000e+02,1.860000000000000000e+02,1.430000000000000000e+02,1.310000000000000000e+02,1.610000000000000000e+02,1.940000000000000000e+02,1.940000000000000000e+02,1.540000000000000000e+02,1.780000000000000000e+02,2.030000000000000000e+02,2.030000000000000000e+02,1.960000000000000000e+02,1.920000000000000000e+02,1.780000000000000000e+02,1.890000000000000000e+02,1.710000000000000000e+02,1.780000000000000000e+02,1.710000000000000000e+02,1.810000000000000000e+02,1.680000000000000000e+02,1.640000000000000000e+02,1.460000000000000000e+02,1.600000000000000000e+02,1.410000000000000000e+02,1.510000000000000000e+02,1.470000000000000000e+02,1.460000000000000000e+02,1.540000000000000000e+02,1.310000000000000000e+02,1.630000000000000000e+02,1.360000000000000000e+02,1.110000000000000000e+02,1.490000000000000000e+02,1.090000000000000000e+02,1.040000000000000000e+02,5.900000000000000000e+01,1.500000000000000000e+01,7.000000000000000000e+00,1.900000000000000000e+01,2.600000000000000000e+01,3.200000000000000000e+01,4.800000000000000000e+01,5.500000000000000000e+01,3.200000000000000000e+01,2.100000000000000000e+01,1.600000000000000000e+01,1.800000000000000000e+01,1.700000000000000000e+01,2.300000000000000000e+01,5.400000000000000000e+01,6.000000000000000000e+01,8.800000000000000000e+01,1.210000000000000000e+02,1.260000000000000000e+02,1.500000000000000000e+02,1.630000000000000000e+02,1.760000000000000000e+02,1.720000000000000000e+02,1.390000000000000000e+02,1.260000000000000000e+02,1.230000000000000000e+02,5.700000000000000000e+01,4.900000000000000000e+01,6.300000000000000000e+01,1.040000000000000000e+02,9.200000000000000000e+01,1.270000000000000000e+02,9.100000000000000000e+01,4.800000000000000000e+01,5.100000000000000000e+01,6.300000000000000000e+01,6.500000000000000000e+01,7.200000000000000000e+01,7.100000000000000000e+01,7.100000000000000000e+01,6.800000000000000000e+01,6.800000000000000000e+01,7.000000000000000000e+01,7.200000000000000000e+01,7.100000000000000000e+01,7.000000000000000000e+01,7.300000000000000000e+01,7.100000000000000000e+01,7.000000000000000000e+01,7.200000000000000000e+01,7.100000000000000000e+01,7.200000000000000000e+01,7.000000000000000000e+01,7.100000000000000000e+01,7.200000000000000000e+01,7.000000000000000000e+01),
(1.490000000000000000e+02,2.000000000000000000e+02,2.070000000000000000e+02,1.990000000000000000e+02,1.900000000000000000e+02,1.750000000000000000e+02,1.570000000000000000e+02,1.410000000000000000e+02,1.420000000000000000e+02,9.100000000000000000e+01,4.100000000000000000e+01,1.400000000000000000e+01,8.000000000000000000e+00,6.000000000000000000e+00,5.000000000000000000e+00,1.500000000000000000e+01,5.500000000000000000e+01,1.520000000000000000e+02,1.650000000000000000e+02,1.610000000000000000e+02,1.500000000000000000e+02,1.770000000000000000e+02,1.400000000000000000e+02,6.200000000000000000e+01,3.000000000000000000e+01,1.200000000000000000e+01,1.600000000000000000e+01,2.400000000000000000e+01,8.000000000000000000e+00,8.000000000000000000e+00,7.000000000000000000e+00,5.800000000000000000e+01,4.900000000000000000e+01,4.800000000000000000e+01,2.200000000000000000e+01,6.600000000000000000e+01,1.010000000000000000e+02,1.240000000000000000e+02,1.200000000000000000e+02,1.290000000000000000e+02,1.540000000000000000e+02,1.910000000000000000e+02,1.590000000000000000e+02,1.420000000000000000e+02,1.640000000000000000e+02,1.940000000000000000e+02,2.030000000000000000e+02,2.000000000000000000e+02,1.890000000000000000e+02,1.740000000000000000e+02,1.770000000000000000e+02,1.940000000000000000e+02,1.760000000000000000e+02,1.970000000000000000e+02,1.760000000000000000e+02,1.880000000000000000e+02,1.800000000000000000e+02,1.640000000000000000e+02,1.710000000000000000e+02,1.610000000000000000e+02,1.560000000000000000e+02,1.480000000000000000e+02,1.760000000000000000e+02,1.380000000000000000e+02,1.430000000000000000e+02,1.620000000000000000e+02,1.600000000000000000e+02,1.480000000000000000e+02,1.280000000000000000e+02,1.290000000000000000e+02,1.330000000000000000e+02,6.900000000000000000e+01,1.800000000000000000e+01,1.800000000000000000e+01,1.800000000000000000e+01,5.300000000000000000e+01,5.300000000000000000e+01,3.600000000000000000e+01,6.400000000000000000e+01,7.200000000000000000e+01,5.400000000000000000e+01,1.600000000000000000e+01,2.000000000000000000e+01,1.700000000000000000e+01,5.300000000000000000e+01,5.200000000000000000e+01,8.900000000000000000e+01,1.060000000000000000e+02,1.220000000000000000e+02,1.480000000000000000e+02,1.380000000000000000e+02,1.380000000000000000e+02,1.190000000000000000e+02,1.410000000000000000e+02,1.530000000000000000e+02,1.410000000000000000e+02,1.040000000000000000e+02,1.070000000000000000e+02,8.000000000000000000e+01,6.800000000000000000e+01,8.800000000000000000e+01,1.090000000000000000e+02,1.190000000000000000e+02,1.210000000000000000e+02,7.300000000000000000e+01,6.300000000000000000e+01,6.900000000000000000e+01,7.700000000000000000e+01,8.900000000000000000e+01,8.900000000000000000e+01,8.600000000000000000e+01,8.900000000000000000e+01,9.000000000000000000e+01,9.100000000000000000e+01,8.700000000000000000e+01,8.700000000000000000e+01,9.200000000000000000e+01,8.700000000000000000e+01,8.700000000000000000e+01,8.600000000000000000e+01,8.800000000000000000e+01,8.700000000000000000e+01,8.400000000000000000e+01,8.600000000000000000e+01,8.200000000000000000e+01,8.600000000000000000e+01,8.100000000000000000e+01,8.500000000000000000e+01),
(1.770000000000000000e+02,2.080000000000000000e+02,2.060000000000000000e+02,1.990000000000000000e+02,1.910000000000000000e+02,1.740000000000000000e+02,1.580000000000000000e+02,1.430000000000000000e+02,1.340000000000000000e+02,1.330000000000000000e+02,1.180000000000000000e+02,3.900000000000000000e+01,2.100000000000000000e+01,7.000000000000000000e+00,5.000000000000000000e+00,1.100000000000000000e+01,1.300000000000000000e+01,2.800000000000000000e+01,7.000000000000000000e+01,1.030000000000000000e+02,1.100000000000000000e+02,1.710000000000000000e+02,1.610000000000000000e+02,8.200000000000000000e+01,3.200000000000000000e+01,2.200000000000000000e+01,2.200000000000000000e+01,2.100000000000000000e+01,1.800000000000000000e+01,1.300000000000000000e+01,2.000000000000000000e+00,4.000000000000000000e+00,1.100000000000000000e+01,1.500000000000000000e+01,2.000000000000000000e+01,3.500000000000000000e+01,5.700000000000000000e+01,8.800000000000000000e+01,1.190000000000000000e+02,1.400000000000000000e+02,1.740000000000000000e+02,1.230000000000000000e+02,1.160000000000000000e+02,1.640000000000000000e+02,1.740000000000000000e+02,1.880000000000000000e+02,1.970000000000000000e+02,1.980000000000000000e+02,1.900000000000000000e+02,1.840000000000000000e+02,1.460000000000000000e+02,1.970000000000000000e+02,1.850000000000000000e+02,2.030000000000000000e+02,1.870000000000000000e+02,1.830000000000000000e+02,1.890000000000000000e+02,1.990000000000000000e+02,1.860000000000000000e+02,1.870000000000000000e+02,1.810000000000000000e+02,1.480000000000000000e+02,1.800000000000000000e+02,1.930000000000000000e+02,1.340000000000000000e+02,1.520000000000000000e+02,1.880000000000000000e+02,1.510000000000000000e+02,1.050000000000000000e+02,8.900000000000000000e+01,9.500000000000000000e+01,3.900000000000000000e+01,1.500000000000000000e+01,2.000000000000000000e+01,6.500000000000000000e+01,4.800000000000000000e+01,3.400000000000000000e+01,1.400000000000000000e+01,2.300000000000000000e+01,5.700000000000000000e+01,3.000000000000000000e+01,3.400000000000000000e+01,2.900000000000000000e+01,3.300000000000000000e+01,6.800000000000000000e+01,1.210000000000000000e+02,1.150000000000000000e+02,1.660000000000000000e+02,1.520000000000000000e+02,1.160000000000000000e+02,1.590000000000000000e+02,1.430000000000000000e+02,1.430000000000000000e+02,8.200000000000000000e+01,6.700000000000000000e+01,8.400000000000000000e+01,1.440000000000000000e+02,1.110000000000000000e+02,5.400000000000000000e+01,5.300000000000000000e+01,6.100000000000000000e+01,8.700000000000000000e+01,1.160000000000000000e+02,1.310000000000000000e+02,7.000000000000000000e+01,4.700000000000000000e+01,7.300000000000000000e+01,9.800000000000000000e+01,9.900000000000000000e+01,9.700000000000000000e+01,1.090000000000000000e+02,1.110000000000000000e+02,9.900000000000000000e+01,1.040000000000000000e+02,1.010000000000000000e+02,1.040000000000000000e+02,1.000000000000000000e+02,1.010000000000000000e+02,9.600000000000000000e+01,9.900000000000000000e+01,1.000000000000000000e+02,9.600000000000000000e+01,9.800000000000000000e+01,9.900000000000000000e+01,9.600000000000000000e+01,9.400000000000000000e+01,9.700000000000000000e+01,9.900000000000000000e+01),
(1.420000000000000000e+02,1.890000000000000000e+02,1.990000000000000000e+02,1.970000000000000000e+02,1.950000000000000000e+02,1.810000000000000000e+02,1.630000000000000000e+02,1.500000000000000000e+02,1.420000000000000000e+02,1.660000000000000000e+02,1.310000000000000000e+02,9.800000000000000000e+01,5.800000000000000000e+01,1.500000000000000000e+01,1.200000000000000000e+01,8.000000000000000000e+00,1.300000000000000000e+01,1.900000000000000000e+01,3.700000000000000000e+01,9.500000000000000000e+01,1.220000000000000000e+02,1.420000000000000000e+02,1.340000000000000000e+02,1.410000000000000000e+02,1.020000000000000000e+02,3.300000000000000000e+01,3.000000000000000000e+01,3.900000000000000000e+01,4.100000000000000000e+01,1.100000000000000000e+01,5.000000000000000000e+00,1.600000000000000000e+01,1.100000000000000000e+01,1.600000000000000000e+01,1.000000000000000000e+01,1.300000000000000000e+01,3.300000000000000000e+01,1.270000000000000000e+02,1.210000000000000000e+02,8.000000000000000000e+01,1.070000000000000000e+02,1.700000000000000000e+02,1.320000000000000000e+02,1.350000000000000000e+02,1.740000000000000000e+02,1.750000000000000000e+02,1.980000000000000000e+02,1.850000000000000000e+02,1.990000000000000000e+02,1.790000000000000000e+02,1.420000000000000000e+02,2.010000000000000000e+02,2.000000000000000000e+02,2.000000000000000000e+02,1.950000000000000000e+02,1.870000000000000000e+02,1.770000000000000000e+02,1.960000000000000000e+02,2.040000000000000000e+02,1.830000000000000000e+02,1.880000000000000000e+02,1.720000000000000000e+02,1.670000000000000000e+02,1.960000000000000000e+02,1.800000000000000000e+02,1.620000000000000000e+02,1.740000000000000000e+02,1.710000000000000000e+02,1.120000000000000000e+02,1.050000000000000000e+02,3.000000000000000000e+01,1.700000000000000000e+01,4.000000000000000000e+01,4.800000000000000000e+01,7.400000000000000000e+01,7.800000000000000000e+01,4.000000000000000000e+01,2.600000000000000000e+01,9.000000000000000000e+00,1.500000000000000000e+01,1.700000000000000000e+01,4.700000000000000000e+01,7.100000000000000000e+01,6.200000000000000000e+01,1.160000000000000000e+02,1.430000000000000000e+02,1.690000000000000000e+02,1.410000000000000000e+02,1.940000000000000000e+02,1.960000000000000000e+02,1.840000000000000000e+02,1.900000000000000000e+02,1.760000000000000000e+02,1.730000000000000000e+02,1.540000000000000000e+02,1.290000000000000000e+02,9.800000000000000000e+01,6.800000000000000000e+01,4.600000000000000000e+01,4.700000000000000000e+01,7.200000000000000000e+01,8.000000000000000000e+01,8.900000000000000000e+01,9.000000000000000000e+01,7.900000000000000000e+01,6.800000000000000000e+01,7.200000000000000000e+01,9.400000000000000000e+01,1.080000000000000000e+02,1.070000000000000000e+02,1.080000000000000000e+02,1.150000000000000000e+02,1.110000000000000000e+02,1.090000000000000000e+02,1.120000000000000000e+02,1.070000000000000000e+02,1.060000000000000000e+02,1.030000000000000000e+02,1.100000000000000000e+02,1.020000000000000000e+02,1.060000000000000000e+02,1.110000000000000000e+02,1.060000000000000000e+02,1.050000000000000000e+02,1.080000000000000000e+02,1.020000000000000000e+02,1.040000000000000000e+02,1.090000000000000000e+02),
(1.370000000000000000e+02,1.890000000000000000e+02,1.980000000000000000e+02,2.010000000000000000e+02,2.030000000000000000e+02,1.980000000000000000e+02,1.840000000000000000e+02,1.590000000000000000e+02,1.690000000000000000e+02,1.810000000000000000e+02,1.560000000000000000e+02,1.620000000000000000e+02,1.500000000000000000e+02,6.600000000000000000e+01,1.700000000000000000e+01,1.900000000000000000e+01,1.000000000000000000e+01,1.500000000000000000e+01,8.000000000000000000e+00,2.600000000000000000e+01,7.000000000000000000e+01,1.200000000000000000e+02,1.400000000000000000e+02,1.350000000000000000e+02,9.500000000000000000e+01,5.800000000000000000e+01,5.100000000000000000e+01,6.300000000000000000e+01,2.500000000000000000e+01,1.300000000000000000e+01,2.300000000000000000e+01,5.100000000000000000e+01,3.000000000000000000e+01,1.200000000000000000e+01,1.300000000000000000e+01,3.400000000000000000e+01,6.000000000000000000e+01,5.300000000000000000e+01,7.400000000000000000e+01,2.900000000000000000e+01,1.090000000000000000e+02,1.570000000000000000e+02,1.330000000000000000e+02,1.540000000000000000e+02,1.900000000000000000e+02,1.650000000000000000e+02,1.880000000000000000e+02,1.890000000000000000e+02,1.810000000000000000e+02,1.610000000000000000e+02,1.250000000000000000e+02,1.810000000000000000e+02,1.990000000000000000e+02,1.990000000000000000e+02,1.970000000000000000e+02,2.040000000000000000e+02,1.700000000000000000e+02,1.950000000000000000e+02,1.960000000000000000e+02,1.840000000000000000e+02,1.790000000000000000e+02,1.960000000000000000e+02,1.520000000000000000e+02,1.530000000000000000e+02,1.990000000000000000e+02,1.580000000000000000e+02,1.440000000000000000e+02,1.730000000000000000e+02,9.200000000000000000e+01,3.700000000000000000e+01,6.600000000000000000e+01,7.200000000000000000e+01,1.120000000000000000e+02,4.100000000000000000e+01,8.600000000000000000e+01,5.600000000000000000e+01,2.400000000000000000e+01,4.300000000000000000e+01,1.900000000000000000e+01,1.500000000000000000e+01,2.400000000000000000e+01,4.700000000000000000e+01,9.600000000000000000e+01,1.390000000000000000e+02,1.110000000000000000e+02,1.500000000000000000e+02,1.670000000000000000e+02,1.980000000000000000e+02,1.780000000000000000e+02,1.400000000000000000e+02,1.260000000000000000e+02,1.510000000000000000e+02,1.480000000000000000e+02,1.240000000000000000e+02,1.590000000000000000e+02,1.450000000000000000e+02,1.030000000000000000e+02,5.800000000000000000e+01,7.200000000000000000e+01,8.400000000000000000e+01,1.060000000000000000e+02,1.440000000000000000e+02,1.110000000000000000e+02,1.380000000000000000e+02,7.600000000000000000e+01,6.400000000000000000e+01,7.700000000000000000e+01,9.300000000000000000e+01,1.010000000000000000e+02,1.070000000000000000e+02,1.100000000000000000e+02,1.180000000000000000e+02,1.140000000000000000e+02,1.180000000000000000e+02,1.190000000000000000e+02,1.130000000000000000e+02,1.130000000000000000e+02,1.110000000000000000e+02,1.120000000000000000e+02,1.090000000000000000e+02,1.110000000000000000e+02,1.100000000000000000e+02,1.080000000000000000e+02,1.080000000000000000e+02,1.070000000000000000e+02,1.090000000000000000e+02,1.080000000000000000e+02,1.070000000000000000e+02),
(1.510000000000000000e+02,1.740000000000000000e+02,1.790000000000000000e+02,1.910000000000000000e+02,1.920000000000000000e+02,1.820000000000000000e+02,1.820000000000000000e+02,1.840000000000000000e+02,2.000000000000000000e+02,2.000000000000000000e+02,1.930000000000000000e+02,1.660000000000000000e+02,1.220000000000000000e+02,8.400000000000000000e+01,5.100000000000000000e+01,2.900000000000000000e+01,1.200000000000000000e+01,4.000000000000000000e+00,1.600000000000000000e+01,5.100000000000000000e+01,3.700000000000000000e+01,8.100000000000000000e+01,1.280000000000000000e+02,1.400000000000000000e+02,1.310000000000000000e+02,1.200000000000000000e+02,6.600000000000000000e+01,4.500000000000000000e+01,5.400000000000000000e+01,3.800000000000000000e+01,8.100000000000000000e+01,7.700000000000000000e+01,6.300000000000000000e+01,5.300000000000000000e+01,1.800000000000000000e+01,3.200000000000000000e+01,3.400000000000000000e+01,4.000000000000000000e+01,1.300000000000000000e+01,5.000000000000000000e+01,6.500000000000000000e+01,9.600000000000000000e+01,1.350000000000000000e+02,1.690000000000000000e+02,1.350000000000000000e+02,1.650000000000000000e+02,1.900000000000000000e+02,1.810000000000000000e+02,1.540000000000000000e+02,1.560000000000000000e+02,1.500000000000000000e+02,1.740000000000000000e+02,2.010000000000000000e+02,1.890000000000000000e+02,1.980000000000000000e+02,2.000000000000000000e+02,1.780000000000000000e+02,1.970000000000000000e+02,1.840000000000000000e+02,1.980000000000000000e+02,1.670000000000000000e+02,1.830000000000000000e+02,1.740000000000000000e+02,1.580000000000000000e+02,1.450000000000000000e+02,1.680000000000000000e+02,9.900000000000000000e+01,1.260000000000000000e+02,8.000000000000000000e+01,8.800000000000000000e+01,1.110000000000000000e+02,1.600000000000000000e+02,7.600000000000000000e+01,7.900000000000000000e+01,1.080000000000000000e+02,3.800000000000000000e+01,1.800000000000000000e+01,1.800000000000000000e+01,2.100000000000000000e+01,2.800000000000000000e+01,3.600000000000000000e+01,6.600000000000000000e+01,1.300000000000000000e+02,1.610000000000000000e+02,1.710000000000000000e+02,1.820000000000000000e+02,1.820000000000000000e+02,1.540000000000000000e+02,9.800000000000000000e+01,1.100000000000000000e+02,8.200000000000000000e+01,1.000000000000000000e+02,1.160000000000000000e+02,8.600000000000000000e+01,3.500000000000000000e+01,5.200000000000000000e+01,3.800000000000000000e+01,4.000000000000000000e+01,4.500000000000000000e+01,9.200000000000000000e+01,1.070000000000000000e+02,1.310000000000000000e+02,1.650000000000000000e+02,1.010000000000000000e+02,5.400000000000000000e+01,5.700000000000000000e+01,8.200000000000000000e+01,9.700000000000000000e+01,1.030000000000000000e+02,1.050000000000000000e+02,1.090000000000000000e+02,1.110000000000000000e+02,1.100000000000000000e+02,1.140000000000000000e+02,1.170000000000000000e+02,1.150000000000000000e+02,1.120000000000000000e+02,1.140000000000000000e+02,1.170000000000000000e+02,1.140000000000000000e+02,1.140000000000000000e+02,1.120000000000000000e+02,1.150000000000000000e+02,1.160000000000000000e+02,1.140000000000000000e+02,1.110000000000000000e+02,1.080000000000000000e+02,1.090000000000000000e+02),
(1.160000000000000000e+02,1.270000000000000000e+02,1.520000000000000000e+02,1.840000000000000000e+02,1.940000000000000000e+02,2.030000000000000000e+02,1.970000000000000000e+02,1.900000000000000000e+02,1.830000000000000000e+02,1.930000000000000000e+02,1.700000000000000000e+02,1.760000000000000000e+02,1.760000000000000000e+02,1.570000000000000000e+02,1.160000000000000000e+02,8.900000000000000000e+01,3.600000000000000000e+01,1.800000000000000000e+01,1.100000000000000000e+01,1.200000000000000000e+01,1.300000000000000000e+01,3.400000000000000000e+01,7.700000000000000000e+01,1.340000000000000000e+02,1.230000000000000000e+02,1.240000000000000000e+02,4.600000000000000000e+01,2.900000000000000000e+01,4.900000000000000000e+01,7.000000000000000000e+01,4.900000000000000000e+01,6.300000000000000000e+01,3.800000000000000000e+01,3.300000000000000000e+01,2.800000000000000000e+01,2.600000000000000000e+01,3.400000000000000000e+01,2.500000000000000000e+01,4.100000000000000000e+01,6.100000000000000000e+01,5.200000000000000000e+01,4.400000000000000000e+01,8.700000000000000000e+01,1.420000000000000000e+02,6.900000000000000000e+01,1.590000000000000000e+02,1.920000000000000000e+02,1.700000000000000000e+02,1.180000000000000000e+02,1.330000000000000000e+02,1.670000000000000000e+02,1.800000000000000000e+02,1.870000000000000000e+02,1.890000000000000000e+02,1.660000000000000000e+02,1.900000000000000000e+02,1.850000000000000000e+02,1.590000000000000000e+02,1.930000000000000000e+02,2.030000000000000000e+02,1.590000000000000000e+02,1.220000000000000000e+02,1.530000000000000000e+02,1.660000000000000000e+02,1.000000000000000000e+02,1.440000000000000000e+02,1.300000000000000000e+02,6.300000000000000000e+01,7.000000000000000000e+01,1.060000000000000000e+02,7.200000000000000000e+01,1.040000000000000000e+02,7.800000000000000000e+01,8.600000000000000000e+01,3.300000000000000000e+01,9.000000000000000000e+00,1.600000000000000000e+01,4.000000000000000000e+01,6.200000000000000000e+01,9.100000000000000000e+01,9.400000000000000000e+01,1.080000000000000000e+02,1.750000000000000000e+02,1.740000000000000000e+02,1.630000000000000000e+02,1.080000000000000000e+02,1.480000000000000000e+02,1.360000000000000000e+02,9.100000000000000000e+01,4.400000000000000000e+01,7.700000000000000000e+01,3.200000000000000000e+01,6.100000000000000000e+01,3.300000000000000000e+01,5.800000000000000000e+01,3.900000000000000000e+01,3.200000000000000000e+01,7.800000000000000000e+01,7.100000000000000000e+01,1.020000000000000000e+02,1.560000000000000000e+02,1.660000000000000000e+02,1.700000000000000000e+02,1.240000000000000000e+02,4.400000000000000000e+01,4.300000000000000000e+01,7.600000000000000000e+01,9.800000000000000000e+01,1.070000000000000000e+02,1.050000000000000000e+02,1.140000000000000000e+02,1.060000000000000000e+02,1.070000000000000000e+02,1.060000000000000000e+02,1.160000000000000000e+02,1.100000000000000000e+02,1.140000000000000000e+02,1.110000000000000000e+02,1.090000000000000000e+02,1.140000000000000000e+02,1.100000000000000000e+02,1.180000000000000000e+02,1.120000000000000000e+02,1.100000000000000000e+02,1.080000000000000000e+02,1.060000000000000000e+02,1.100000000000000000e+02,1.100000000000000000e+02),
(1.400000000000000000e+02,1.800000000000000000e+02,1.870000000000000000e+02,1.860000000000000000e+02,1.840000000000000000e+02,1.840000000000000000e+02,1.900000000000000000e+02,1.880000000000000000e+02,1.990000000000000000e+02,1.980000000000000000e+02,1.760000000000000000e+02,1.400000000000000000e+02,1.960000000000000000e+02,1.970000000000000000e+02,1.860000000000000000e+02,1.640000000000000000e+02,1.030000000000000000e+02,6.400000000000000000e+01,2.500000000000000000e+01,9.000000000000000000e+00,7.000000000000000000e+00,4.000000000000000000e+00,1.100000000000000000e+01,7.000000000000000000e+01,1.300000000000000000e+02,1.550000000000000000e+02,7.300000000000000000e+01,6.100000000000000000e+01,4.800000000000000000e+01,2.700000000000000000e+01,7.200000000000000000e+01,7.400000000000000000e+01,4.700000000000000000e+01,6.500000000000000000e+01,8.000000000000000000e+01,6.900000000000000000e+01,8.000000000000000000e+01,4.600000000000000000e+01,3.100000000000000000e+01,2.500000000000000000e+01,7.400000000000000000e+01,6.800000000000000000e+01,7.200000000000000000e+01,1.060000000000000000e+02,4.500000000000000000e+01,1.080000000000000000e+02,1.480000000000000000e+02,1.220000000000000000e+02,6.000000000000000000e+01,1.110000000000000000e+02,1.820000000000000000e+02,1.900000000000000000e+02,1.960000000000000000e+02,1.890000000000000000e+02,1.660000000000000000e+02,1.650000000000000000e+02,1.900000000000000000e+02,1.700000000000000000e+02,1.690000000000000000e+02,1.480000000000000000e+02,1.420000000000000000e+02,1.260000000000000000e+02,9.600000000000000000e+01,1.720000000000000000e+02,1.180000000000000000e+02,5.500000000000000000e+01,1.420000000000000000e+02,8.400000000000000000e+01,9.500000000000000000e+01,1.060000000000000000e+02,1.190000000000000000e+02,8.300000000000000000e+01,5.300000000000000000e+01,3.500000000000000000e+01,1.700000000000000000e+01,1.100000000000000000e+01,2.900000000000000000e+01,6.900000000000000000e+01,1.040000000000000000e+02,1.000000000000000000e+02,1.250000000000000000e+02,1.320000000000000000e+02,1.670000000000000000e+02,1.820000000000000000e+02,1.310000000000000000e+02,1.620000000000000000e+02,1.330000000000000000e+02,1.030000000000000000e+02,6.200000000000000000e+01,4.800000000000000000e+01,1.800000000000000000e+01,4.600000000000000000e+01,2.600000000000000000e+01,2.400000000000000000e+01,4.200000000000000000e+01,6.900000000000000000e+01,5.500000000000000000e+01,1.190000000000000000e+02,1.500000000000000000e+02,1.360000000000000000e+02,1.130000000000000000e+02,1.530000000000000000e+02,1.540000000000000000e+02,1.160000000000000000e+02,9.000000000000000000e+01,5.900000000000000000e+01,7.300000000000000000e+01,8.600000000000000000e+01,9.800000000000000000e+01,1.020000000000000000e+02,1.080000000000000000e+02,1.090000000000000000e+02,1.040000000000000000e+02,1.060000000000000000e+02,1.050000000000000000e+02,1.060000000000000000e+02,1.080000000000000000e+02,1.080000000000000000e+02,1.080000000000000000e+02,1.120000000000000000e+02,1.090000000000000000e+02,1.110000000000000000e+02,1.100000000000000000e+02,1.090000000000000000e+02,1.060000000000000000e+02,1.050000000000000000e+02,1.110000000000000000e+02,1.070000000000000000e+02),
(1.450000000000000000e+02,1.010000000000000000e+02,9.700000000000000000e+01,1.530000000000000000e+02,1.610000000000000000e+02,1.680000000000000000e+02,1.650000000000000000e+02,1.700000000000000000e+02,1.910000000000000000e+02,1.920000000000000000e+02,1.800000000000000000e+02,1.680000000000000000e+02,1.820000000000000000e+02,1.950000000000000000e+02,1.780000000000000000e+02,1.490000000000000000e+02,1.400000000000000000e+02,9.000000000000000000e+01,4.300000000000000000e+01,1.700000000000000000e+01,9.000000000000000000e+00,3.000000000000000000e+00,4.000000000000000000e+00,3.600000000000000000e+01,1.010000000000000000e+02,1.220000000000000000e+02,1.430000000000000000e+02,8.000000000000000000e+01,6.600000000000000000e+01,7.800000000000000000e+01,3.500000000000000000e+01,6.800000000000000000e+01,9.200000000000000000e+01,1.130000000000000000e+02,1.290000000000000000e+02,6.300000000000000000e+01,7.700000000000000000e+01,4.100000000000000000e+01,5.300000000000000000e+01,4.400000000000000000e+01,5.500000000000000000e+01,4.600000000000000000e+01,9.100000000000000000e+01,5.500000000000000000e+01,6.000000000000000000e+01,1.250000000000000000e+02,1.030000000000000000e+02,1.090000000000000000e+02,2.900000000000000000e+01,1.150000000000000000e+02,1.890000000000000000e+02,1.590000000000000000e+02,1.760000000000000000e+02,1.860000000000000000e+02,1.510000000000000000e+02,1.400000000000000000e+02,1.920000000000000000e+02,2.080000000000000000e+02,1.710000000000000000e+02,1.040000000000000000e+02,1.410000000000000000e+02,1.580000000000000000e+02,1.170000000000000000e+02,9.500000000000000000e+01,8.700000000000000000e+01,6.700000000000000000e+01,9.000000000000000000e+01,1.190000000000000000e+02,1.560000000000000000e+02,1.460000000000000000e+02,3.700000000000000000e+01,8.900000000000000000e+01,2.400000000000000000e+01,3.100000000000000000e+01,2.900000000000000000e+01,4.000000000000000000e+01,9.700000000000000000e+01,6.800000000000000000e+01,1.070000000000000000e+02,1.280000000000000000e+02,1.800000000000000000e+02,1.300000000000000000e+02,1.640000000000000000e+02,1.600000000000000000e+02,1.720000000000000000e+02,1.420000000000000000e+02,1.550000000000000000e+02,1.330000000000000000e+02,1.020000000000000000e+02,9.300000000000000000e+01,9.200000000000000000e+01,3.500000000000000000e+01,8.000000000000000000e+00,1.900000000000000000e+01,3.600000000000000000e+01,3.700000000000000000e+01,1.260000000000000000e+02,1.620000000000000000e+02,1.750000000000000000e+02,1.720000000000000000e+02,1.560000000000000000e+02,1.570000000000000000e+02,1.750000000000000000e+02,1.160000000000000000e+02,2.900000000000000000e+01,3.000000000000000000e+01,6.400000000000000000e+01,7.900000000000000000e+01,9.300000000000000000e+01,9.800000000000000000e+01,1.010000000000000000e+02,1.010000000000000000e+02,9.700000000000000000e+01,1.060000000000000000e+02,1.000000000000000000e+02,1.060000000000000000e+02,1.020000000000000000e+02,9.900000000000000000e+01,1.030000000000000000e+02,1.050000000000000000e+02,1.060000000000000000e+02,1.050000000000000000e+02,1.050000000000000000e+02,1.030000000000000000e+02,1.040000000000000000e+02,1.020000000000000000e+02,1.040000000000000000e+02,1.030000000000000000e+02),
(1.600000000000000000e+02,1.540000000000000000e+02,1.790000000000000000e+02,1.970000000000000000e+02,2.020000000000000000e+02,1.940000000000000000e+02,1.840000000000000000e+02,1.890000000000000000e+02,1.780000000000000000e+02,1.910000000000000000e+02,1.840000000000000000e+02,1.660000000000000000e+02,1.650000000000000000e+02,1.940000000000000000e+02,1.970000000000000000e+02,1.840000000000000000e+02,1.580000000000000000e+02,1.470000000000000000e+02,1.220000000000000000e+02,3.900000000000000000e+01,1.900000000000000000e+01,8.000000000000000000e+00,8.000000000000000000e+00,2.700000000000000000e+01,6.700000000000000000e+01,1.350000000000000000e+02,1.100000000000000000e+02,8.300000000000000000e+01,5.900000000000000000e+01,5.300000000000000000e+01,8.300000000000000000e+01,1.150000000000000000e+02,1.290000000000000000e+02,1.820000000000000000e+02,1.050000000000000000e+02,1.110000000000000000e+02,9.500000000000000000e+01,8.700000000000000000e+01,8.400000000000000000e+01,8.000000000000000000e+01,8.500000000000000000e+01,6.100000000000000000e+01,7.300000000000000000e+01,5.200000000000000000e+01,9.300000000000000000e+01,1.350000000000000000e+02,9.100000000000000000e+01,1.000000000000000000e+02,4.700000000000000000e+01,9.300000000000000000e+01,1.340000000000000000e+02,1.750000000000000000e+02,1.510000000000000000e+02,1.590000000000000000e+02,1.230000000000000000e+02,1.360000000000000000e+02,1.330000000000000000e+02,2.020000000000000000e+02,1.740000000000000000e+02,1.150000000000000000e+02,1.320000000000000000e+02,1.760000000000000000e+02,1.390000000000000000e+02,1.290000000000000000e+02,7.200000000000000000e+01,7.200000000000000000e+01,1.230000000000000000e+02,1.540000000000000000e+02,2.000000000000000000e+02,1.570000000000000000e+02,1.700000000000000000e+01,2.800000000000000000e+01,4.200000000000000000e+01,2.900000000000000000e+01,7.000000000000000000e+01,7.500000000000000000e+01,1.350000000000000000e+02,1.380000000000000000e+02,1.620000000000000000e+02,1.390000000000000000e+02,1.580000000000000000e+02,1.520000000000000000e+02,1.610000000000000000e+02,1.650000000000000000e+02,1.440000000000000000e+02,1.360000000000000000e+02,1.000000000000000000e+02,1.510000000000000000e+02,8.000000000000000000e+01,2.600000000000000000e+01,3.600000000000000000e+01,3.000000000000000000e+01,2.100000000000000000e+01,3.300000000000000000e+01,9.500000000000000000e+01,9.900000000000000000e+01,1.200000000000000000e+02,1.950000000000000000e+02,1.940000000000000000e+02,1.590000000000000000e+02,1.500000000000000000e+02,1.490000000000000000e+02,1.380000000000000000e+02,7.700000000000000000e+01,3.100000000000000000e+01,2.800000000000000000e+01,5.400000000000000000e+01,7.900000000000000000e+01,8.300000000000000000e+01,8.900000000000000000e+01,9.300000000000000000e+01,9.700000000000000000e+01,9.500000000000000000e+01,9.700000000000000000e+01,9.800000000000000000e+01,1.000000000000000000e+02,9.600000000000000000e+01,1.020000000000000000e+02,9.900000000000000000e+01,9.700000000000000000e+01,1.010000000000000000e+02,1.080000000000000000e+02,9.700000000000000000e+01,9.600000000000000000e+01,1.020000000000000000e+02,1.010000000000000000e+02,9.800000000000000000e+01,9.900000000000000000e+01),
(1.530000000000000000e+02,1.480000000000000000e+02,1.530000000000000000e+02,1.740000000000000000e+02,1.870000000000000000e+02,1.860000000000000000e+02,1.950000000000000000e+02,1.930000000000000000e+02,1.810000000000000000e+02,1.790000000000000000e+02,1.750000000000000000e+02,1.540000000000000000e+02,1.760000000000000000e+02,1.800000000000000000e+02,1.800000000000000000e+02,1.800000000000000000e+02,1.480000000000000000e+02,1.640000000000000000e+02,1.730000000000000000e+02,1.060000000000000000e+02,9.000000000000000000e+01,7.100000000000000000e+01,1.600000000000000000e+01,7.000000000000000000e+00,2.400000000000000000e+01,8.800000000000000000e+01,1.560000000000000000e+02,1.240000000000000000e+02,8.800000000000000000e+01,5.200000000000000000e+01,2.700000000000000000e+01,5.000000000000000000e+01,9.300000000000000000e+01,1.220000000000000000e+02,1.410000000000000000e+02,8.800000000000000000e+01,1.000000000000000000e+02,1.120000000000000000e+02,1.430000000000000000e+02,7.900000000000000000e+01,1.220000000000000000e+02,1.440000000000000000e+02,7.600000000000000000e+01,5.700000000000000000e+01,8.300000000000000000e+01,1.130000000000000000e+02,9.700000000000000000e+01,8.100000000000000000e+01,6.200000000000000000e+01,1.110000000000000000e+02,7.600000000000000000e+01,1.500000000000000000e+02,1.230000000000000000e+02,7.400000000000000000e+01,6.900000000000000000e+01,1.430000000000000000e+02,1.770000000000000000e+02,1.050000000000000000e+02,1.610000000000000000e+02,1.310000000000000000e+02,1.100000000000000000e+02,1.110000000000000000e+02,1.020000000000000000e+02,9.500000000000000000e+01,6.600000000000000000e+01,9.900000000000000000e+01,1.380000000000000000e+02,1.420000000000000000e+02,1.370000000000000000e+02,9.400000000000000000e+01,3.300000000000000000e+01,2.300000000000000000e+01,6.000000000000000000e+01,1.240000000000000000e+02,9.400000000000000000e+01,9.300000000000000000e+01,9.200000000000000000e+01,1.570000000000000000e+02,1.550000000000000000e+02,1.800000000000000000e+02,1.350000000000000000e+02,1.750000000000000000e+02,7.400000000000000000e+01,1.680000000000000000e+02,1.150000000000000000e+02,7.300000000000000000e+01,6.100000000000000000e+01,5.100000000000000000e+01,4.300000000000000000e+01,3.400000000000000000e+01,3.000000000000000000e+01,2.700000000000000000e+01,4.300000000000000000e+01,8.000000000000000000e+01,1.060000000000000000e+02,1.300000000000000000e+02,1.490000000000000000e+02,1.440000000000000000e+02,1.560000000000000000e+02,1.780000000000000000e+02,1.940000000000000000e+02,1.890000000000000000e+02,1.170000000000000000e+02,3.900000000000000000e+01,1.300000000000000000e+01,1.500000000000000000e+01,4.100000000000000000e+01,7.900000000000000000e+01,8.900000000000000000e+01,8.800000000000000000e+01,9.200000000000000000e+01,9.100000000000000000e+01,9.000000000000000000e+01,9.400000000000000000e+01,9.300000000000000000e+01,9.400000000000000000e+01,9.100000000000000000e+01,9.500000000000000000e+01,9.300000000000000000e+01,9.400000000000000000e+01,9.500000000000000000e+01,9.400000000000000000e+01,9.600000000000000000e+01,9.700000000000000000e+01,9.900000000000000000e+01,9.700000000000000000e+01,9.800000000000000000e+01,9.900000000000000000e+01),
(1.570000000000000000e+02,1.560000000000000000e+02,1.220000000000000000e+02,1.340000000000000000e+02,9.900000000000000000e+01,9.600000000000000000e+01,1.480000000000000000e+02,1.470000000000000000e+02,1.450000000000000000e+02,1.630000000000000000e+02,1.640000000000000000e+02,1.520000000000000000e+02,1.710000000000000000e+02,1.790000000000000000e+02,1.820000000000000000e+02,1.560000000000000000e+02,1.250000000000000000e+02,1.450000000000000000e+02,1.500000000000000000e+02,1.630000000000000000e+02,1.500000000000000000e+02,9.000000000000000000e+01,3.400000000000000000e+01,1.400000000000000000e+01,1.400000000000000000e+01,5.400000000000000000e+01,1.470000000000000000e+02,1.740000000000000000e+02,1.500000000000000000e+02,1.100000000000000000e+02,5.400000000000000000e+01,5.800000000000000000e+01,9.700000000000000000e+01,8.200000000000000000e+01,6.500000000000000000e+01,1.120000000000000000e+02,1.670000000000000000e+02,1.480000000000000000e+02,1.180000000000000000e+02,8.400000000000000000e+01,1.050000000000000000e+02,1.280000000000000000e+02,1.200000000000000000e+02,1.180000000000000000e+02,9.800000000000000000e+01,9.300000000000000000e+01,1.210000000000000000e+02,1.450000000000000000e+02,1.030000000000000000e+02,1.090000000000000000e+02,1.100000000000000000e+02,1.070000000000000000e+02,1.500000000000000000e+02,1.110000000000000000e+02,1.020000000000000000e+02,8.800000000000000000e+01,1.520000000000000000e+02,1.090000000000000000e+02,8.900000000000000000e+01,1.350000000000000000e+02,1.120000000000000000e+02,8.900000000000000000e+01,8.400000000000000000e+01,1.040000000000000000e+02,1.220000000000000000e+02,1.120000000000000000e+02,1.400000000000000000e+02,1.520000000000000000e+02,9.900000000000000000e+01,3.400000000000000000e+01,8.400000000000000000e+01,8.100000000000000000e+01,6.800000000000000000e+01,1.190000000000000000e+02,1.140000000000000000e+02,1.150000000000000000e+02,8.600000000000000000e+01,9.800000000000000000e+01,1.810000000000000000e+02,1.490000000000000000e+02,1.140000000000000000e+02,1.010000000000000000e+02,1.190000000000000000e+02,7.500000000000000000e+01,9.100000000000000000e+01,5.400000000000000000e+01,8.500000000000000000e+01,2.200000000000000000e+01,3.100000000000000000e+01,1.900000000000000000e+01,2.100000000000000000e+01,4.400000000000000000e+01,7.600000000000000000e+01,1.440000000000000000e+02,1.450000000000000000e+02,1.080000000000000000e+02,1.150000000000000000e+02,1.680000000000000000e+02,1.610000000000000000e+02,1.400000000000000000e+02,1.490000000000000000e+02,1.580000000000000000e+02,1.490000000000000000e+02,4.000000000000000000e+01,1.400000000000000000e+01,1.400000000000000000e+01,2.200000000000000000e+01,6.300000000000000000e+01,8.400000000000000000e+01,8.700000000000000000e+01,8.900000000000000000e+01,9.300000000000000000e+01,8.800000000000000000e+01,9.300000000000000000e+01,8.700000000000000000e+01,8.900000000000000000e+01,9.100000000000000000e+01,9.200000000000000000e+01,8.900000000000000000e+01,9.300000000000000000e+01,9.200000000000000000e+01,9.100000000000000000e+01,9.200000000000000000e+01,9.600000000000000000e+01,9.600000000000000000e+01,9.700000000000000000e+01,9.600000000000000000e+01,9.200000000000000000e+01),
(1.640000000000000000e+02,1.390000000000000000e+02,9.100000000000000000e+01,5.900000000000000000e+01,6.100000000000000000e+01,6.100000000000000000e+01,9.000000000000000000e+01,8.400000000000000000e+01,1.390000000000000000e+02,1.660000000000000000e+02,1.750000000000000000e+02,1.770000000000000000e+02,1.790000000000000000e+02,1.480000000000000000e+02,1.480000000000000000e+02,1.440000000000000000e+02,1.260000000000000000e+02,1.150000000000000000e+02,1.380000000000000000e+02,1.630000000000000000e+02,1.520000000000000000e+02,1.200000000000000000e+02,7.900000000000000000e+01,7.100000000000000000e+01,2.100000000000000000e+01,1.300000000000000000e+01,4.300000000000000000e+01,6.700000000000000000e+01,1.600000000000000000e+02,1.090000000000000000e+02,1.040000000000000000e+02,9.600000000000000000e+01,3.900000000000000000e+01,1.900000000000000000e+01,6.900000000000000000e+01,1.530000000000000000e+02,1.270000000000000000e+02,1.840000000000000000e+02,1.270000000000000000e+02,1.270000000000000000e+02,1.350000000000000000e+02,1.330000000000000000e+02,1.550000000000000000e+02,1.580000000000000000e+02,1.360000000000000000e+02,1.160000000000000000e+02,1.690000000000000000e+02,1.340000000000000000e+02,1.370000000000000000e+02,1.240000000000000000e+02,1.200000000000000000e+02,1.200000000000000000e+02,1.370000000000000000e+02,1.530000000000000000e+02,8.000000000000000000e+01,8.700000000000000000e+01,1.220000000000000000e+02,8.100000000000000000e+01,6.800000000000000000e+01,1.020000000000000000e+02,8.500000000000000000e+01,9.300000000000000000e+01,1.090000000000000000e+02,1.150000000000000000e+02,1.520000000000000000e+02,1.180000000000000000e+02,1.330000000000000000e+02,1.070000000000000000e+02,4.000000000000000000e+01,7.900000000000000000e+01,1.260000000000000000e+02,1.510000000000000000e+02,1.620000000000000000e+02,1.210000000000000000e+02,9.900000000000000000e+01,6.700000000000000000e+01,1.260000000000000000e+02,7.300000000000000000e+01,1.290000000000000000e+02,1.140000000000000000e+02,9.000000000000000000e+01,1.180000000000000000e+02,1.070000000000000000e+02,1.500000000000000000e+01,2.600000000000000000e+01,3.900000000000000000e+01,6.600000000000000000e+01,3.700000000000000000e+01,1.100000000000000000e+01,4.500000000000000000e+01,8.500000000000000000e+01,6.900000000000000000e+01,8.500000000000000000e+01,1.240000000000000000e+02,1.640000000000000000e+02,1.160000000000000000e+02,1.490000000000000000e+02,1.390000000000000000e+02,1.490000000000000000e+02,1.390000000000000000e+02,1.410000000000000000e+02,4.500000000000000000e+01,3.000000000000000000e+01,2.700000000000000000e+01,1.800000000000000000e+01,2.200000000000000000e+01,2.200000000000000000e+01,4.900000000000000000e+01,7.900000000000000000e+01,8.500000000000000000e+01,8.500000000000000000e+01,8.500000000000000000e+01,9.000000000000000000e+01,8.600000000000000000e+01,8.900000000000000000e+01,9.200000000000000000e+01,8.300000000000000000e+01,8.800000000000000000e+01,8.900000000000000000e+01,9.200000000000000000e+01,9.000000000000000000e+01,8.800000000000000000e+01,9.000000000000000000e+01,8.800000000000000000e+01,9.700000000000000000e+01,9.200000000000000000e+01,9.800000000000000000e+01,9.700000000000000000e+01),
(1.620000000000000000e+02,1.520000000000000000e+02,1.180000000000000000e+02,1.210000000000000000e+02,1.170000000000000000e+02,9.400000000000000000e+01,8.500000000000000000e+01,1.030000000000000000e+02,1.610000000000000000e+02,1.680000000000000000e+02,1.770000000000000000e+02,1.940000000000000000e+02,1.840000000000000000e+02,1.800000000000000000e+02,1.720000000000000000e+02,1.630000000000000000e+02,1.750000000000000000e+02,1.790000000000000000e+02,1.560000000000000000e+02,1.750000000000000000e+02,1.880000000000000000e+02,1.580000000000000000e+02,1.300000000000000000e+02,8.700000000000000000e+01,4.100000000000000000e+01,1.400000000000000000e+01,7.000000000000000000e+00,2.800000000000000000e+01,1.230000000000000000e+02,1.190000000000000000e+02,1.200000000000000000e+02,1.010000000000000000e+02,6.000000000000000000e+01,6.600000000000000000e+01,8.100000000000000000e+01,1.010000000000000000e+02,1.420000000000000000e+02,1.550000000000000000e+02,1.570000000000000000e+02,1.780000000000000000e+02,1.470000000000000000e+02,1.890000000000000000e+02,1.530000000000000000e+02,1.730000000000000000e+02,1.520000000000000000e+02,1.730000000000000000e+02,1.580000000000000000e+02,1.090000000000000000e+02,1.510000000000000000e+02,1.770000000000000000e+02,1.730000000000000000e+02,1.380000000000000000e+02,1.550000000000000000e+02,1.580000000000000000e+02,1.160000000000000000e+02,1.340000000000000000e+02,1.290000000000000000e+02,1.060000000000000000e+02,1.010000000000000000e+02,1.420000000000000000e+02,1.530000000000000000e+02,1.150000000000000000e+02,1.430000000000000000e+02,1.600000000000000000e+02,2.020000000000000000e+02,1.600000000000000000e+02,1.530000000000000000e+02,3.200000000000000000e+01,2.700000000000000000e+01,1.580000000000000000e+02,1.250000000000000000e+02,1.210000000000000000e+02,1.480000000000000000e+02,1.950000000000000000e+02,1.250000000000000000e+02,1.260000000000000000e+02,1.500000000000000000e+02,1.100000000000000000e+02,1.230000000000000000e+02,1.420000000000000000e+02,1.390000000000000000e+02,8.600000000000000000e+01,5.400000000000000000e+01,1.400000000000000000e+01,4.000000000000000000e+00,8.000000000000000000e+00,1.800000000000000000e+01,2.300000000000000000e+01,3.200000000000000000e+01,4.800000000000000000e+01,8.200000000000000000e+01,1.590000000000000000e+02,1.890000000000000000e+02,1.640000000000000000e+02,1.510000000000000000e+02,1.460000000000000000e+02,1.520000000000000000e+02,1.760000000000000000e+02,1.630000000000000000e+02,1.220000000000000000e+02,9.200000000000000000e+01,4.700000000000000000e+01,1.000000000000000000e+01,9.000000000000000000e+00,1.000000000000000000e+01,1.800000000000000000e+01,2.200000000000000000e+01,4.200000000000000000e+01,7.700000000000000000e+01,8.800000000000000000e+01,8.900000000000000000e+01,9.200000000000000000e+01,9.000000000000000000e+01,8.300000000000000000e+01,8.600000000000000000e+01,8.600000000000000000e+01,8.800000000000000000e+01,8.600000000000000000e+01,9.100000000000000000e+01,8.700000000000000000e+01,9.000000000000000000e+01,8.800000000000000000e+01,9.200000000000000000e+01,9.000000000000000000e+01,9.100000000000000000e+01,9.200000000000000000e+01,9.500000000000000000e+01,9.400000000000000000e+01),
(1.570000000000000000e+02,1.600000000000000000e+02,1.660000000000000000e+02,1.690000000000000000e+02,1.380000000000000000e+02,1.160000000000000000e+02,1.410000000000000000e+02,1.760000000000000000e+02,1.740000000000000000e+02,1.720000000000000000e+02,1.780000000000000000e+02,1.810000000000000000e+02,1.870000000000000000e+02,1.760000000000000000e+02,1.830000000000000000e+02,1.910000000000000000e+02,1.650000000000000000e+02,1.400000000000000000e+02,1.510000000000000000e+02,1.430000000000000000e+02,1.520000000000000000e+02,1.880000000000000000e+02,1.600000000000000000e+02,1.660000000000000000e+02,8.700000000000000000e+01,5.700000000000000000e+01,1.100000000000000000e+01,1.800000000000000000e+01,6.800000000000000000e+01,1.550000000000000000e+02,1.200000000000000000e+02,9.700000000000000000e+01,9.000000000000000000e+01,6.100000000000000000e+01,5.700000000000000000e+01,7.900000000000000000e+01,9.900000000000000000e+01,1.540000000000000000e+02,1.930000000000000000e+02,1.380000000000000000e+02,2.020000000000000000e+02,1.940000000000000000e+02,1.900000000000000000e+02,1.690000000000000000e+02,1.920000000000000000e+02,1.790000000000000000e+02,1.810000000000000000e+02,1.820000000000000000e+02,1.560000000000000000e+02,1.930000000000000000e+02,1.610000000000000000e+02,1.810000000000000000e+02,1.680000000000000000e+02,1.900000000000000000e+02,1.600000000000000000e+02,1.280000000000000000e+02,1.400000000000000000e+02,1.590000000000000000e+02,1.570000000000000000e+02,1.840000000000000000e+02,1.760000000000000000e+02,1.720000000000000000e+02,1.810000000000000000e+02,2.110000000000000000e+02,2.090000000000000000e+02,1.590000000000000000e+02,1.380000000000000000e+02,9.500000000000000000e+01,5.800000000000000000e+01,1.620000000000000000e+02,1.290000000000000000e+02,1.580000000000000000e+02,1.260000000000000000e+02,1.920000000000000000e+02,1.210000000000000000e+02,9.800000000000000000e+01,1.590000000000000000e+02,8.500000000000000000e+01,2.900000000000000000e+01,5.600000000000000000e+01,1.270000000000000000e+02,3.000000000000000000e+01,3.400000000000000000e+01,2.500000000000000000e+01,1.500000000000000000e+01,1.700000000000000000e+01,1.700000000000000000e+01,2.700000000000000000e+01,8.800000000000000000e+01,1.040000000000000000e+02,1.440000000000000000e+02,1.560000000000000000e+02,1.890000000000000000e+02,2.040000000000000000e+02,1.780000000000000000e+02,1.720000000000000000e+02,1.480000000000000000e+02,1.920000000000000000e+02,1.610000000000000000e+02,1.190000000000000000e+02,5.800000000000000000e+01,3.500000000000000000e+01,1.200000000000000000e+01,9.000000000000000000e+00,1.000000000000000000e+01,1.500000000000000000e+01,2.700000000000000000e+01,3.800000000000000000e+01,7.200000000000000000e+01,8.600000000000000000e+01,9.200000000000000000e+01,9.100000000000000000e+01,8.600000000000000000e+01,8.800000000000000000e+01,8.700000000000000000e+01,8.700000000000000000e+01,9.000000000000000000e+01,8.600000000000000000e+01,9.100000000000000000e+01,8.700000000000000000e+01,8.700000000000000000e+01,8.800000000000000000e+01,8.800000000000000000e+01,8.800000000000000000e+01,9.400000000000000000e+01,9.000000000000000000e+01,9.400000000000000000e+01,9.400000000000000000e+01),
(1.900000000000000000e+02,1.920000000000000000e+02,1.910000000000000000e+02,1.620000000000000000e+02,1.410000000000000000e+02,1.120000000000000000e+02,1.140000000000000000e+02,1.620000000000000000e+02,1.700000000000000000e+02,1.790000000000000000e+02,1.670000000000000000e+02,1.590000000000000000e+02,1.590000000000000000e+02,1.510000000000000000e+02,1.880000000000000000e+02,1.890000000000000000e+02,1.670000000000000000e+02,1.550000000000000000e+02,1.570000000000000000e+02,1.650000000000000000e+02,1.520000000000000000e+02,1.410000000000000000e+02,1.500000000000000000e+02,1.490000000000000000e+02,1.320000000000000000e+02,1.180000000000000000e+02,4.200000000000000000e+01,8.000000000000000000e+00,1.200000000000000000e+01,5.300000000000000000e+01,1.360000000000000000e+02,1.490000000000000000e+02,1.210000000000000000e+02,2.400000000000000000e+01,9.900000000000000000e+01,1.090000000000000000e+02,8.400000000000000000e+01,1.250000000000000000e+02,1.110000000000000000e+02,1.660000000000000000e+02,1.830000000000000000e+02,1.880000000000000000e+02,1.620000000000000000e+02,1.770000000000000000e+02,1.780000000000000000e+02,1.380000000000000000e+02,1.670000000000000000e+02,1.890000000000000000e+02,1.770000000000000000e+02,1.870000000000000000e+02,1.860000000000000000e+02,1.910000000000000000e+02,1.950000000000000000e+02,2.040000000000000000e+02,1.930000000000000000e+02,1.890000000000000000e+02,2.010000000000000000e+02,1.970000000000000000e+02,1.830000000000000000e+02,1.890000000000000000e+02,2.010000000000000000e+02,1.980000000000000000e+02,1.800000000000000000e+02,2.030000000000000000e+02,2.030000000000000000e+02,1.620000000000000000e+02,1.590000000000000000e+02,1.150000000000000000e+02,7.400000000000000000e+01,1.390000000000000000e+02,1.310000000000000000e+02,1.300000000000000000e+02,1.440000000000000000e+02,1.030000000000000000e+02,4.000000000000000000e+01,5.900000000000000000e+01,3.500000000000000000e+01,1.200000000000000000e+01,2.600000000000000000e+01,1.800000000000000000e+01,1.200000000000000000e+01,4.000000000000000000e+01,3.500000000000000000e+01,1.200000000000000000e+01,4.400000000000000000e+01,3.200000000000000000e+01,7.900000000000000000e+01,4.500000000000000000e+01,1.160000000000000000e+02,1.650000000000000000e+02,1.840000000000000000e+02,1.620000000000000000e+02,1.660000000000000000e+02,1.980000000000000000e+02,1.760000000000000000e+02,1.770000000000000000e+02,1.380000000000000000e+02,8.700000000000000000e+01,1.250000000000000000e+02,1.510000000000000000e+02,7.300000000000000000e+01,1.700000000000000000e+01,1.400000000000000000e+01,1.400000000000000000e+01,8.000000000000000000e+00,2.300000000000000000e+01,3.000000000000000000e+01,2.900000000000000000e+01,6.200000000000000000e+01,8.500000000000000000e+01,8.900000000000000000e+01,9.300000000000000000e+01,9.000000000000000000e+01,8.800000000000000000e+01,9.000000000000000000e+01,9.000000000000000000e+01,8.700000000000000000e+01,8.600000000000000000e+01,8.900000000000000000e+01,8.600000000000000000e+01,8.700000000000000000e+01,9.000000000000000000e+01,9.100000000000000000e+01,9.400000000000000000e+01,9.500000000000000000e+01,9.800000000000000000e+01,9.700000000000000000e+01,9.700000000000000000e+01));
     END PROCESS tb;
  END;
